module switch(
    input [67:0]bits0,
    input [67:0]bits1,
    input [67:0]bits2,
    input [67:0]bits3,
    input [67:0]bits4,
    input [67:0]bits5,
    input [67:0]bits6,
    input [67:0]bits7,
    input [67:0]bits8,
    input [67:0]bits9,
    input [67:0]bits10,
    input [67:0]bits11,
    input [67:0]bits12,
    input [67:0]bits13,
    input [67:0]bits14,
    input [67:0]bits15,
    input [67:0]bits16,
    output [16:0]exbits0,
    output [16:0]exbits1,
    output [16:0]exbits2,
    output [16:0]exbits3,
    output [16:0]exbits4,
    output [16:0]exbits5,
    output [16:0]exbits6,
    output [16:0]exbits7,
    output [16:0]exbits8,
    output [16:0]exbits9,
    output [16:0]exbits10,
    output [16:0]exbits11,
    output [16:0]exbits12,
    output [16:0]exbits13,
    output [16:0]exbits14,
    output [16:0]exbits15,
    output [16:0]exbits16,
    output [16:0]exbits17,
    output [16:0]exbits18,
    output [16:0]exbits19,
    output [16:0]exbits20,
    output [16:0]exbits21,
    output [16:0]exbits22,
    output [16:0]exbits23,
    output [16:0]exbits24,
    output [16:0]exbits25,
    output [16:0]exbits26,
    output [16:0]exbits27,
    output [16:0]exbits28,
    output [16:0]exbits29,
    output [16:0]exbits30,
    output [16:0]exbits31,
    output [16:0]exbits32,
    output [16:0]exbits33,
    output [16:0]exbits34,
    output [16:0]exbits35,
    output [16:0]exbits36,
    output [16:0]exbits37,
    output [16:0]exbits38,
    output [16:0]exbits39,
    output [16:0]exbits40,
    output [16:0]exbits41,
    output [16:0]exbits42,
    output [16:0]exbits43,
    output [16:0]exbits44,
    output [16:0]exbits45,
    output [16:0]exbits46,
    output [16:0]exbits47,
    output [16:0]exbits48,
    output [16:0]exbits49,
    output [16:0]exbits50,
    output [16:0]exbits51,
    output [16:0]exbits52,
    output [16:0]exbits53,
    output [16:0]exbits54,
    output [16:0]exbits55,
    output [16:0]exbits56,
    output [16:0]exbits57,
    output [16:0]exbits58,
    output [16:0]exbits59,
    output [16:0]exbits60,
    output [16:0]exbits61,
    output [16:0]exbits62,
    output [16:0]exbits63,
    output [16:0]exbits64,
    output [16:0]exbits65,
    output [16:0]exbits66,
    output [16:0]exbits67
);
assign exbits0 = {
bits0[0],
bits1[0],
bits2[0],
bits3[0],
bits4[0],
bits5[0],
bits6[0],
bits7[0],
bits8[0],
bits9[0],
bits10[0],
bits11[0],
bits12[0],
bits13[0],
bits14[0],
bits15[0],
bits16[0]};

assign exbits1 = {
bits0[1],
bits1[1],
bits2[1],
bits3[1],
bits4[1],
bits5[1],
bits6[1],
bits7[1],
bits8[1],
bits9[1],
bits10[1],
bits11[1],
bits12[1],
bits13[1],
bits14[1],
bits15[1],
bits16[1]};

assign exbits2 = {
bits0[2],
bits1[2],
bits2[2],
bits3[2],
bits4[2],
bits5[2],
bits6[2],
bits7[2],
bits8[2],
bits9[2],
bits10[2],
bits11[2],
bits12[2],
bits13[2],
bits14[2],
bits15[2],
bits16[2]};

assign exbits3 = {
bits0[3],
bits1[3],
bits2[3],
bits3[3],
bits4[3],
bits5[3],
bits6[3],
bits7[3],
bits8[3],
bits9[3],
bits10[3],
bits11[3],
bits12[3],
bits13[3],
bits14[3],
bits15[3],
bits16[3]};

assign exbits4 = {
bits0[4],
bits1[4],
bits2[4],
bits3[4],
bits4[4],
bits5[4],
bits6[4],
bits7[4],
bits8[4],
bits9[4],
bits10[4],
bits11[4],
bits12[4],
bits13[4],
bits14[4],
bits15[4],
bits16[4]};

assign exbits5 = {
bits0[5],
bits1[5],
bits2[5],
bits3[5],
bits4[5],
bits5[5],
bits6[5],
bits7[5],
bits8[5],
bits9[5],
bits10[5],
bits11[5],
bits12[5],
bits13[5],
bits14[5],
bits15[5],
bits16[5]};

assign exbits6 = {
bits0[6],
bits1[6],
bits2[6],
bits3[6],
bits4[6],
bits5[6],
bits6[6],
bits7[6],
bits8[6],
bits9[6],
bits10[6],
bits11[6],
bits12[6],
bits13[6],
bits14[6],
bits15[6],
bits16[6]};

assign exbits7 = {
bits0[7],
bits1[7],
bits2[7],
bits3[7],
bits4[7],
bits5[7],
bits6[7],
bits7[7],
bits8[7],
bits9[7],
bits10[7],
bits11[7],
bits12[7],
bits13[7],
bits14[7],
bits15[7],
bits16[7]};

assign exbits8 = {
bits0[8],
bits1[8],
bits2[8],
bits3[8],
bits4[8],
bits5[8],
bits6[8],
bits7[8],
bits8[8],
bits9[8],
bits10[8],
bits11[8],
bits12[8],
bits13[8],
bits14[8],
bits15[8],
bits16[8]};

assign exbits9 = {
bits0[9],
bits1[9],
bits2[9],
bits3[9],
bits4[9],
bits5[9],
bits6[9],
bits7[9],
bits8[9],
bits9[9],
bits10[9],
bits11[9],
bits12[9],
bits13[9],
bits14[9],
bits15[9],
bits16[9]};

assign exbits10 = {
bits0[10],
bits1[10],
bits2[10],
bits3[10],
bits4[10],
bits5[10],
bits6[10],
bits7[10],
bits8[10],
bits9[10],
bits10[10],
bits11[10],
bits12[10],
bits13[10],
bits14[10],
bits15[10],
bits16[10]};

assign exbits11 = {
bits0[11],
bits1[11],
bits2[11],
bits3[11],
bits4[11],
bits5[11],
bits6[11],
bits7[11],
bits8[11],
bits9[11],
bits10[11],
bits11[11],
bits12[11],
bits13[11],
bits14[11],
bits15[11],
bits16[11]};

assign exbits12 = {
bits0[12],
bits1[12],
bits2[12],
bits3[12],
bits4[12],
bits5[12],
bits6[12],
bits7[12],
bits8[12],
bits9[12],
bits10[12],
bits11[12],
bits12[12],
bits13[12],
bits14[12],
bits15[12],
bits16[12]};

assign exbits13 = {
bits0[13],
bits1[13],
bits2[13],
bits3[13],
bits4[13],
bits5[13],
bits6[13],
bits7[13],
bits8[13],
bits9[13],
bits10[13],
bits11[13],
bits12[13],
bits13[13],
bits14[13],
bits15[13],
bits16[13]};

assign exbits14 = {
bits0[14],
bits1[14],
bits2[14],
bits3[14],
bits4[14],
bits5[14],
bits6[14],
bits7[14],
bits8[14],
bits9[14],
bits10[14],
bits11[14],
bits12[14],
bits13[14],
bits14[14],
bits15[14],
bits16[14]};

assign exbits15 = {
bits0[15],
bits1[15],
bits2[15],
bits3[15],
bits4[15],
bits5[15],
bits6[15],
bits7[15],
bits8[15],
bits9[15],
bits10[15],
bits11[15],
bits12[15],
bits13[15],
bits14[15],
bits15[15],
bits16[15]};

assign exbits16 = {
bits0[16],
bits1[16],
bits2[16],
bits3[16],
bits4[16],
bits5[16],
bits6[16],
bits7[16],
bits8[16],
bits9[16],
bits10[16],
bits11[16],
bits12[16],
bits13[16],
bits14[16],
bits15[16],
bits16[16]};

assign exbits17 = {
bits0[17],
bits1[17],
bits2[17],
bits3[17],
bits4[17],
bits5[17],
bits6[17],
bits7[17],
bits8[17],
bits9[17],
bits10[17],
bits11[17],
bits12[17],
bits13[17],
bits14[17],
bits15[17],
bits16[17]};

assign exbits18 = {
bits0[18],
bits1[18],
bits2[18],
bits3[18],
bits4[18],
bits5[18],
bits6[18],
bits7[18],
bits8[18],
bits9[18],
bits10[18],
bits11[18],
bits12[18],
bits13[18],
bits14[18],
bits15[18],
bits16[18]};

assign exbits19 = {
bits0[19],
bits1[19],
bits2[19],
bits3[19],
bits4[19],
bits5[19],
bits6[19],
bits7[19],
bits8[19],
bits9[19],
bits10[19],
bits11[19],
bits12[19],
bits13[19],
bits14[19],
bits15[19],
bits16[19]};

assign exbits20 = {
bits0[20],
bits1[20],
bits2[20],
bits3[20],
bits4[20],
bits5[20],
bits6[20],
bits7[20],
bits8[20],
bits9[20],
bits10[20],
bits11[20],
bits12[20],
bits13[20],
bits14[20],
bits15[20],
bits16[20]};

assign exbits21 = {
bits0[21],
bits1[21],
bits2[21],
bits3[21],
bits4[21],
bits5[21],
bits6[21],
bits7[21],
bits8[21],
bits9[21],
bits10[21],
bits11[21],
bits12[21],
bits13[21],
bits14[21],
bits15[21],
bits16[21]};

assign exbits22 = {
bits0[22],
bits1[22],
bits2[22],
bits3[22],
bits4[22],
bits5[22],
bits6[22],
bits7[22],
bits8[22],
bits9[22],
bits10[22],
bits11[22],
bits12[22],
bits13[22],
bits14[22],
bits15[22],
bits16[22]};

assign exbits23 = {
bits0[23],
bits1[23],
bits2[23],
bits3[23],
bits4[23],
bits5[23],
bits6[23],
bits7[23],
bits8[23],
bits9[23],
bits10[23],
bits11[23],
bits12[23],
bits13[23],
bits14[23],
bits15[23],
bits16[23]};

assign exbits24 = {
bits0[24],
bits1[24],
bits2[24],
bits3[24],
bits4[24],
bits5[24],
bits6[24],
bits7[24],
bits8[24],
bits9[24],
bits10[24],
bits11[24],
bits12[24],
bits13[24],
bits14[24],
bits15[24],
bits16[24]};

assign exbits25 = {
bits0[25],
bits1[25],
bits2[25],
bits3[25],
bits4[25],
bits5[25],
bits6[25],
bits7[25],
bits8[25],
bits9[25],
bits10[25],
bits11[25],
bits12[25],
bits13[25],
bits14[25],
bits15[25],
bits16[25]};

assign exbits26 = {
bits0[26],
bits1[26],
bits2[26],
bits3[26],
bits4[26],
bits5[26],
bits6[26],
bits7[26],
bits8[26],
bits9[26],
bits10[26],
bits11[26],
bits12[26],
bits13[26],
bits14[26],
bits15[26],
bits16[26]};

assign exbits27 = {
bits0[27],
bits1[27],
bits2[27],
bits3[27],
bits4[27],
bits5[27],
bits6[27],
bits7[27],
bits8[27],
bits9[27],
bits10[27],
bits11[27],
bits12[27],
bits13[27],
bits14[27],
bits15[27],
bits16[27]};

assign exbits28 = {
bits0[28],
bits1[28],
bits2[28],
bits3[28],
bits4[28],
bits5[28],
bits6[28],
bits7[28],
bits8[28],
bits9[28],
bits10[28],
bits11[28],
bits12[28],
bits13[28],
bits14[28],
bits15[28],
bits16[28]};

assign exbits29 = {
bits0[29],
bits1[29],
bits2[29],
bits3[29],
bits4[29],
bits5[29],
bits6[29],
bits7[29],
bits8[29],
bits9[29],
bits10[29],
bits11[29],
bits12[29],
bits13[29],
bits14[29],
bits15[29],
bits16[29]};

assign exbits30 = {
bits0[30],
bits1[30],
bits2[30],
bits3[30],
bits4[30],
bits5[30],
bits6[30],
bits7[30],
bits8[30],
bits9[30],
bits10[30],
bits11[30],
bits12[30],
bits13[30],
bits14[30],
bits15[30],
bits16[30]};

assign exbits31 = {
bits0[31],
bits1[31],
bits2[31],
bits3[31],
bits4[31],
bits5[31],
bits6[31],
bits7[31],
bits8[31],
bits9[31],
bits10[31],
bits11[31],
bits12[31],
bits13[31],
bits14[31],
bits15[31],
bits16[31]};

assign exbits32 = {
bits0[32],
bits1[32],
bits2[32],
bits3[32],
bits4[32],
bits5[32],
bits6[32],
bits7[32],
bits8[32],
bits9[32],
bits10[32],
bits11[32],
bits12[32],
bits13[32],
bits14[32],
bits15[32],
bits16[32]};

assign exbits33 = {
bits0[33],
bits1[33],
bits2[33],
bits3[33],
bits4[33],
bits5[33],
bits6[33],
bits7[33],
bits8[33],
bits9[33],
bits10[33],
bits11[33],
bits12[33],
bits13[33],
bits14[33],
bits15[33],
bits16[33]};

assign exbits34 = {
bits0[34],
bits1[34],
bits2[34],
bits3[34],
bits4[34],
bits5[34],
bits6[34],
bits7[34],
bits8[34],
bits9[34],
bits10[34],
bits11[34],
bits12[34],
bits13[34],
bits14[34],
bits15[34],
bits16[34]};

assign exbits35 = {
bits0[35],
bits1[35],
bits2[35],
bits3[35],
bits4[35],
bits5[35],
bits6[35],
bits7[35],
bits8[35],
bits9[35],
bits10[35],
bits11[35],
bits12[35],
bits13[35],
bits14[35],
bits15[35],
bits16[35]};

assign exbits36 = {
bits0[36],
bits1[36],
bits2[36],
bits3[36],
bits4[36],
bits5[36],
bits6[36],
bits7[36],
bits8[36],
bits9[36],
bits10[36],
bits11[36],
bits12[36],
bits13[36],
bits14[36],
bits15[36],
bits16[36]};

assign exbits37 = {
bits0[37],
bits1[37],
bits2[37],
bits3[37],
bits4[37],
bits5[37],
bits6[37],
bits7[37],
bits8[37],
bits9[37],
bits10[37],
bits11[37],
bits12[37],
bits13[37],
bits14[37],
bits15[37],
bits16[37]};

assign exbits38 = {
bits0[38],
bits1[38],
bits2[38],
bits3[38],
bits4[38],
bits5[38],
bits6[38],
bits7[38],
bits8[38],
bits9[38],
bits10[38],
bits11[38],
bits12[38],
bits13[38],
bits14[38],
bits15[38],
bits16[38]};

assign exbits39 = {
bits0[39],
bits1[39],
bits2[39],
bits3[39],
bits4[39],
bits5[39],
bits6[39],
bits7[39],
bits8[39],
bits9[39],
bits10[39],
bits11[39],
bits12[39],
bits13[39],
bits14[39],
bits15[39],
bits16[39]};

assign exbits40 = {
bits0[40],
bits1[40],
bits2[40],
bits3[40],
bits4[40],
bits5[40],
bits6[40],
bits7[40],
bits8[40],
bits9[40],
bits10[40],
bits11[40],
bits12[40],
bits13[40],
bits14[40],
bits15[40],
bits16[40]};

assign exbits41 = {
bits0[41],
bits1[41],
bits2[41],
bits3[41],
bits4[41],
bits5[41],
bits6[41],
bits7[41],
bits8[41],
bits9[41],
bits10[41],
bits11[41],
bits12[41],
bits13[41],
bits14[41],
bits15[41],
bits16[41]};

assign exbits42 = {
bits0[42],
bits1[42],
bits2[42],
bits3[42],
bits4[42],
bits5[42],
bits6[42],
bits7[42],
bits8[42],
bits9[42],
bits10[42],
bits11[42],
bits12[42],
bits13[42],
bits14[42],
bits15[42],
bits16[42]};

assign exbits43 = {
bits0[43],
bits1[43],
bits2[43],
bits3[43],
bits4[43],
bits5[43],
bits6[43],
bits7[43],
bits8[43],
bits9[43],
bits10[43],
bits11[43],
bits12[43],
bits13[43],
bits14[43],
bits15[43],
bits16[43]};

assign exbits44 = {
bits0[44],
bits1[44],
bits2[44],
bits3[44],
bits4[44],
bits5[44],
bits6[44],
bits7[44],
bits8[44],
bits9[44],
bits10[44],
bits11[44],
bits12[44],
bits13[44],
bits14[44],
bits15[44],
bits16[44]};

assign exbits45 = {
bits0[45],
bits1[45],
bits2[45],
bits3[45],
bits4[45],
bits5[45],
bits6[45],
bits7[45],
bits8[45],
bits9[45],
bits10[45],
bits11[45],
bits12[45],
bits13[45],
bits14[45],
bits15[45],
bits16[45]};

assign exbits46 = {
bits0[46],
bits1[46],
bits2[46],
bits3[46],
bits4[46],
bits5[46],
bits6[46],
bits7[46],
bits8[46],
bits9[46],
bits10[46],
bits11[46],
bits12[46],
bits13[46],
bits14[46],
bits15[46],
bits16[46]};

assign exbits47 = {
bits0[47],
bits1[47],
bits2[47],
bits3[47],
bits4[47],
bits5[47],
bits6[47],
bits7[47],
bits8[47],
bits9[47],
bits10[47],
bits11[47],
bits12[47],
bits13[47],
bits14[47],
bits15[47],
bits16[47]};

assign exbits48 = {
bits0[48],
bits1[48],
bits2[48],
bits3[48],
bits4[48],
bits5[48],
bits6[48],
bits7[48],
bits8[48],
bits9[48],
bits10[48],
bits11[48],
bits12[48],
bits13[48],
bits14[48],
bits15[48],
bits16[48]};

assign exbits49 = {
bits0[49],
bits1[49],
bits2[49],
bits3[49],
bits4[49],
bits5[49],
bits6[49],
bits7[49],
bits8[49],
bits9[49],
bits10[49],
bits11[49],
bits12[49],
bits13[49],
bits14[49],
bits15[49],
bits16[49]};

assign exbits50 = {
bits0[50],
bits1[50],
bits2[50],
bits3[50],
bits4[50],
bits5[50],
bits6[50],
bits7[50],
bits8[50],
bits9[50],
bits10[50],
bits11[50],
bits12[50],
bits13[50],
bits14[50],
bits15[50],
bits16[50]};

assign exbits51 = {
bits0[51],
bits1[51],
bits2[51],
bits3[51],
bits4[51],
bits5[51],
bits6[51],
bits7[51],
bits8[51],
bits9[51],
bits10[51],
bits11[51],
bits12[51],
bits13[51],
bits14[51],
bits15[51],
bits16[51]};

assign exbits52 = {
bits0[52],
bits1[52],
bits2[52],
bits3[52],
bits4[52],
bits5[52],
bits6[52],
bits7[52],
bits8[52],
bits9[52],
bits10[52],
bits11[52],
bits12[52],
bits13[52],
bits14[52],
bits15[52],
bits16[52]};

assign exbits53 = {
bits0[53],
bits1[53],
bits2[53],
bits3[53],
bits4[53],
bits5[53],
bits6[53],
bits7[53],
bits8[53],
bits9[53],
bits10[53],
bits11[53],
bits12[53],
bits13[53],
bits14[53],
bits15[53],
bits16[53]};

assign exbits54 = {
bits0[54],
bits1[54],
bits2[54],
bits3[54],
bits4[54],
bits5[54],
bits6[54],
bits7[54],
bits8[54],
bits9[54],
bits10[54],
bits11[54],
bits12[54],
bits13[54],
bits14[54],
bits15[54],
bits16[54]};

assign exbits55 = {
bits0[55],
bits1[55],
bits2[55],
bits3[55],
bits4[55],
bits5[55],
bits6[55],
bits7[55],
bits8[55],
bits9[55],
bits10[55],
bits11[55],
bits12[55],
bits13[55],
bits14[55],
bits15[55],
bits16[55]};

assign exbits56 = {
bits0[56],
bits1[56],
bits2[56],
bits3[56],
bits4[56],
bits5[56],
bits6[56],
bits7[56],
bits8[56],
bits9[56],
bits10[56],
bits11[56],
bits12[56],
bits13[56],
bits14[56],
bits15[56],
bits16[56]};

assign exbits57 = {
bits0[57],
bits1[57],
bits2[57],
bits3[57],
bits4[57],
bits5[57],
bits6[57],
bits7[57],
bits8[57],
bits9[57],
bits10[57],
bits11[57],
bits12[57],
bits13[57],
bits14[57],
bits15[57],
bits16[57]};

assign exbits58 = {
bits0[58],
bits1[58],
bits2[58],
bits3[58],
bits4[58],
bits5[58],
bits6[58],
bits7[58],
bits8[58],
bits9[58],
bits10[58],
bits11[58],
bits12[58],
bits13[58],
bits14[58],
bits15[58],
bits16[58]};

assign exbits59 = {
bits0[59],
bits1[59],
bits2[59],
bits3[59],
bits4[59],
bits5[59],
bits6[59],
bits7[59],
bits8[59],
bits9[59],
bits10[59],
bits11[59],
bits12[59],
bits13[59],
bits14[59],
bits15[59],
bits16[59]};

assign exbits60 = {
bits0[60],
bits1[60],
bits2[60],
bits3[60],
bits4[60],
bits5[60],
bits6[60],
bits7[60],
bits8[60],
bits9[60],
bits10[60],
bits11[60],
bits12[60],
bits13[60],
bits14[60],
bits15[60],
bits16[60]};

assign exbits61 = {
bits0[61],
bits1[61],
bits2[61],
bits3[61],
bits4[61],
bits5[61],
bits6[61],
bits7[61],
bits8[61],
bits9[61],
bits10[61],
bits11[61],
bits12[61],
bits13[61],
bits14[61],
bits15[61],
bits16[61]};

assign exbits62 = {
bits0[62],
bits1[62],
bits2[62],
bits3[62],
bits4[62],
bits5[62],
bits6[62],
bits7[62],
bits8[62],
bits9[62],
bits10[62],
bits11[62],
bits12[62],
bits13[62],
bits14[62],
bits15[62],
bits16[62]};

assign exbits63 = {
bits0[63],
bits1[63],
bits2[63],
bits3[63],
bits4[63],
bits5[63],
bits6[63],
bits7[63],
bits8[63],
bits9[63],
bits10[63],
bits11[63],
bits12[63],
bits13[63],
bits14[63],
bits15[63],
bits16[63]};

assign exbits64 = {
bits0[64],
bits1[64],
bits2[64],
bits3[64],
bits4[64],
bits5[64],
bits6[64],
bits7[64],
bits8[64],
bits9[64],
bits10[64],
bits11[64],
bits12[64],
bits13[64],
bits14[64],
bits15[64],
bits16[64]};

assign exbits65 = {
bits0[65],
bits1[65],
bits2[65],
bits3[65],
bits4[65],
bits5[65],
bits6[65],
bits7[65],
bits8[65],
bits9[65],
bits10[65],
bits11[65],
bits12[65],
bits13[65],
bits14[65],
bits15[65],
bits16[65]};

assign exbits66 = {
bits0[66],
bits1[66],
bits2[66],
bits3[66],
bits4[66],
bits5[66],
bits6[66],
bits7[66],
bits8[66],
bits9[66],
bits10[66],
bits11[66],
bits12[66],
bits13[66],
bits14[66],
bits15[66],
bits16[66]};

assign exbits67 = {
bits0[67],
bits1[67],
bits2[67],
bits3[67],
bits4[67],
bits5[67],
bits6[67],
bits7[67],
bits8[67],
bits9[67],
bits10[67],
bits11[67],
bits12[67],
bits13[67],
bits14[67],
bits15[67],
bits16[67]};


endmodule