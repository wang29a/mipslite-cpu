
module controller_uint(
    input wire [5:0]op;
    output RegDst,
    output Branch,
    output MemRead,
    output MemtoReg,
    output [1:0] ALUOp,
    output Memwrite,
    output ALUsrc,
    output RegWrite
);

endmodule