`include "head.v"
`include "part_product-template.v"
`include "special_part_product.v"
`include "get_c.v"
`include "switch.v"
`include "walloc_17bits-template.v"
`include "cla_68bits.v"
module multiplier(
    input sign,
    input [31:0] _X,
    input [31:0] _Y,
    output  [63:0] res,
    output reg [67:0] extend_X
);
wire [67:0] part_p [0:16];
// reg [11:0] extend_X;
reg [67:0] move_ex[0:16];
reg [34:0] Y;
// wire [1:0]C[0:16];
wire [67:0]C;
integer i, j;
always @(*) 
begin
    if(sign == 1'b0)
    begin
        extend_X = {36'b0, _X};
        Y = {2'b0, _Y, 1'b0};
    end
    else
    begin
      extend_X = {{36{_X[31]}}, _X};
      Y = {{2{_Y[31]}}, _Y, 1'b0};
    end  
    for(i = 0; i < 17; i = i + 1)
        move_ex[i] = extend_X << (2 *( i));

    // res = 0;
    // for(i = 0; i < 17; i = i + 1)
    // begin
    //     res = res + part_p[i];
    //     res = res + (C[i] << (i * 2));
    // end
    
end
s_part_product sp0000(move_ex[0][0:0], Y[2:0], part_p[0][0]);
part_product p0001(move_ex[0][1:0], Y[2:0], part_p[0][1]);
part_product p0002(move_ex[0][2:1], Y[2:0], part_p[0][2]);
part_product p0003(move_ex[0][3:2], Y[2:0], part_p[0][3]);
part_product p0004(move_ex[0][4:3], Y[2:0], part_p[0][4]);
part_product p0005(move_ex[0][5:4], Y[2:0], part_p[0][5]);
part_product p0006(move_ex[0][6:5], Y[2:0], part_p[0][6]);
part_product p0007(move_ex[0][7:6], Y[2:0], part_p[0][7]);
part_product p0008(move_ex[0][8:7], Y[2:0], part_p[0][8]);
part_product p0009(move_ex[0][9:8], Y[2:0], part_p[0][9]);
part_product p0010(move_ex[0][10:9], Y[2:0], part_p[0][10]);
part_product p0011(move_ex[0][11:10], Y[2:0], part_p[0][11]);
part_product p0012(move_ex[0][12:11], Y[2:0], part_p[0][12]);
part_product p0013(move_ex[0][13:12], Y[2:0], part_p[0][13]);
part_product p0014(move_ex[0][14:13], Y[2:0], part_p[0][14]);
part_product p0015(move_ex[0][15:14], Y[2:0], part_p[0][15]);
part_product p0016(move_ex[0][16:15], Y[2:0], part_p[0][16]);
part_product p0017(move_ex[0][17:16], Y[2:0], part_p[0][17]);
part_product p0018(move_ex[0][18:17], Y[2:0], part_p[0][18]);
part_product p0019(move_ex[0][19:18], Y[2:0], part_p[0][19]);
part_product p0020(move_ex[0][20:19], Y[2:0], part_p[0][20]);
part_product p0021(move_ex[0][21:20], Y[2:0], part_p[0][21]);
part_product p0022(move_ex[0][22:21], Y[2:0], part_p[0][22]);
part_product p0023(move_ex[0][23:22], Y[2:0], part_p[0][23]);
part_product p0024(move_ex[0][24:23], Y[2:0], part_p[0][24]);
part_product p0025(move_ex[0][25:24], Y[2:0], part_p[0][25]);
part_product p0026(move_ex[0][26:25], Y[2:0], part_p[0][26]);
part_product p0027(move_ex[0][27:26], Y[2:0], part_p[0][27]);
part_product p0028(move_ex[0][28:27], Y[2:0], part_p[0][28]);
part_product p0029(move_ex[0][29:28], Y[2:0], part_p[0][29]);
part_product p0030(move_ex[0][30:29], Y[2:0], part_p[0][30]);
part_product p0031(move_ex[0][31:30], Y[2:0], part_p[0][31]);
part_product p0032(move_ex[0][32:31], Y[2:0], part_p[0][32]);
part_product p0033(move_ex[0][33:32], Y[2:0], part_p[0][33]);
part_product p0034(move_ex[0][34:33], Y[2:0], part_p[0][34]);
part_product p0035(move_ex[0][35:34], Y[2:0], part_p[0][35]);
part_product p0036(move_ex[0][36:35], Y[2:0], part_p[0][36]);
part_product p0037(move_ex[0][37:36], Y[2:0], part_p[0][37]);
part_product p0038(move_ex[0][38:37], Y[2:0], part_p[0][38]);
part_product p0039(move_ex[0][39:38], Y[2:0], part_p[0][39]);
part_product p0040(move_ex[0][40:39], Y[2:0], part_p[0][40]);
part_product p0041(move_ex[0][41:40], Y[2:0], part_p[0][41]);
part_product p0042(move_ex[0][42:41], Y[2:0], part_p[0][42]);
part_product p0043(move_ex[0][43:42], Y[2:0], part_p[0][43]);
part_product p0044(move_ex[0][44:43], Y[2:0], part_p[0][44]);
part_product p0045(move_ex[0][45:44], Y[2:0], part_p[0][45]);
part_product p0046(move_ex[0][46:45], Y[2:0], part_p[0][46]);
part_product p0047(move_ex[0][47:46], Y[2:0], part_p[0][47]);
part_product p0048(move_ex[0][48:47], Y[2:0], part_p[0][48]);
part_product p0049(move_ex[0][49:48], Y[2:0], part_p[0][49]);
part_product p0050(move_ex[0][50:49], Y[2:0], part_p[0][50]);
part_product p0051(move_ex[0][51:50], Y[2:0], part_p[0][51]);
part_product p0052(move_ex[0][52:51], Y[2:0], part_p[0][52]);
part_product p0053(move_ex[0][53:52], Y[2:0], part_p[0][53]);
part_product p0054(move_ex[0][54:53], Y[2:0], part_p[0][54]);
part_product p0055(move_ex[0][55:54], Y[2:0], part_p[0][55]);
part_product p0056(move_ex[0][56:55], Y[2:0], part_p[0][56]);
part_product p0057(move_ex[0][57:56], Y[2:0], part_p[0][57]);
part_product p0058(move_ex[0][58:57], Y[2:0], part_p[0][58]);
part_product p0059(move_ex[0][59:58], Y[2:0], part_p[0][59]);
part_product p0060(move_ex[0][60:59], Y[2:0], part_p[0][60]);
part_product p0061(move_ex[0][61:60], Y[2:0], part_p[0][61]);
part_product p0062(move_ex[0][62:61], Y[2:0], part_p[0][62]);
part_product p0063(move_ex[0][63:62], Y[2:0], part_p[0][63]);
part_product p0064(move_ex[0][64:63], Y[2:0], part_p[0][64]);
part_product p0065(move_ex[0][65:64], Y[2:0], part_p[0][65]);
part_product p0066(move_ex[0][66:65], Y[2:0], part_p[0][66]);
part_product p0067(move_ex[0][67:66], Y[2:0], part_p[0][67]);
get_c getc0(Y[2:0], C[1:0]);

assign part_p[1][0] = 0;
assign part_p[1][1] = 0;
s_part_product sp0102(move_ex[1][2:2], Y[4:2], part_p[1][2]);
part_product p0103(move_ex[1][3:2], Y[4:2], part_p[1][3]);
part_product p0104(move_ex[1][4:3], Y[4:2], part_p[1][4]);
part_product p0105(move_ex[1][5:4], Y[4:2], part_p[1][5]);
part_product p0106(move_ex[1][6:5], Y[4:2], part_p[1][6]);
part_product p0107(move_ex[1][7:6], Y[4:2], part_p[1][7]);
part_product p0108(move_ex[1][8:7], Y[4:2], part_p[1][8]);
part_product p0109(move_ex[1][9:8], Y[4:2], part_p[1][9]);
part_product p0110(move_ex[1][10:9], Y[4:2], part_p[1][10]);
part_product p0111(move_ex[1][11:10], Y[4:2], part_p[1][11]);
part_product p0112(move_ex[1][12:11], Y[4:2], part_p[1][12]);
part_product p0113(move_ex[1][13:12], Y[4:2], part_p[1][13]);
part_product p0114(move_ex[1][14:13], Y[4:2], part_p[1][14]);
part_product p0115(move_ex[1][15:14], Y[4:2], part_p[1][15]);
part_product p0116(move_ex[1][16:15], Y[4:2], part_p[1][16]);
part_product p0117(move_ex[1][17:16], Y[4:2], part_p[1][17]);
part_product p0118(move_ex[1][18:17], Y[4:2], part_p[1][18]);
part_product p0119(move_ex[1][19:18], Y[4:2], part_p[1][19]);
part_product p0120(move_ex[1][20:19], Y[4:2], part_p[1][20]);
part_product p0121(move_ex[1][21:20], Y[4:2], part_p[1][21]);
part_product p0122(move_ex[1][22:21], Y[4:2], part_p[1][22]);
part_product p0123(move_ex[1][23:22], Y[4:2], part_p[1][23]);
part_product p0124(move_ex[1][24:23], Y[4:2], part_p[1][24]);
part_product p0125(move_ex[1][25:24], Y[4:2], part_p[1][25]);
part_product p0126(move_ex[1][26:25], Y[4:2], part_p[1][26]);
part_product p0127(move_ex[1][27:26], Y[4:2], part_p[1][27]);
part_product p0128(move_ex[1][28:27], Y[4:2], part_p[1][28]);
part_product p0129(move_ex[1][29:28], Y[4:2], part_p[1][29]);
part_product p0130(move_ex[1][30:29], Y[4:2], part_p[1][30]);
part_product p0131(move_ex[1][31:30], Y[4:2], part_p[1][31]);
part_product p0132(move_ex[1][32:31], Y[4:2], part_p[1][32]);
part_product p0133(move_ex[1][33:32], Y[4:2], part_p[1][33]);
part_product p0134(move_ex[1][34:33], Y[4:2], part_p[1][34]);
part_product p0135(move_ex[1][35:34], Y[4:2], part_p[1][35]);
part_product p0136(move_ex[1][36:35], Y[4:2], part_p[1][36]);
part_product p0137(move_ex[1][37:36], Y[4:2], part_p[1][37]);
part_product p0138(move_ex[1][38:37], Y[4:2], part_p[1][38]);
part_product p0139(move_ex[1][39:38], Y[4:2], part_p[1][39]);
part_product p0140(move_ex[1][40:39], Y[4:2], part_p[1][40]);
part_product p0141(move_ex[1][41:40], Y[4:2], part_p[1][41]);
part_product p0142(move_ex[1][42:41], Y[4:2], part_p[1][42]);
part_product p0143(move_ex[1][43:42], Y[4:2], part_p[1][43]);
part_product p0144(move_ex[1][44:43], Y[4:2], part_p[1][44]);
part_product p0145(move_ex[1][45:44], Y[4:2], part_p[1][45]);
part_product p0146(move_ex[1][46:45], Y[4:2], part_p[1][46]);
part_product p0147(move_ex[1][47:46], Y[4:2], part_p[1][47]);
part_product p0148(move_ex[1][48:47], Y[4:2], part_p[1][48]);
part_product p0149(move_ex[1][49:48], Y[4:2], part_p[1][49]);
part_product p0150(move_ex[1][50:49], Y[4:2], part_p[1][50]);
part_product p0151(move_ex[1][51:50], Y[4:2], part_p[1][51]);
part_product p0152(move_ex[1][52:51], Y[4:2], part_p[1][52]);
part_product p0153(move_ex[1][53:52], Y[4:2], part_p[1][53]);
part_product p0154(move_ex[1][54:53], Y[4:2], part_p[1][54]);
part_product p0155(move_ex[1][55:54], Y[4:2], part_p[1][55]);
part_product p0156(move_ex[1][56:55], Y[4:2], part_p[1][56]);
part_product p0157(move_ex[1][57:56], Y[4:2], part_p[1][57]);
part_product p0158(move_ex[1][58:57], Y[4:2], part_p[1][58]);
part_product p0159(move_ex[1][59:58], Y[4:2], part_p[1][59]);
part_product p0160(move_ex[1][60:59], Y[4:2], part_p[1][60]);
part_product p0161(move_ex[1][61:60], Y[4:2], part_p[1][61]);
part_product p0162(move_ex[1][62:61], Y[4:2], part_p[1][62]);
part_product p0163(move_ex[1][63:62], Y[4:2], part_p[1][63]);
part_product p0164(move_ex[1][64:63], Y[4:2], part_p[1][64]);
part_product p0165(move_ex[1][65:64], Y[4:2], part_p[1][65]);
part_product p0166(move_ex[1][66:65], Y[4:2], part_p[1][66]);
part_product p0167(move_ex[1][67:66], Y[4:2], part_p[1][67]);
get_c getc1(Y[4:2], C[3:2]);

assign part_p[2][0] = 0;
assign part_p[2][1] = 0;
assign part_p[2][2] = 0;
assign part_p[2][3] = 0;
s_part_product sp0204(move_ex[2][4:4], Y[6:4], part_p[2][4]);
part_product p0205(move_ex[2][5:4], Y[6:4], part_p[2][5]);
part_product p0206(move_ex[2][6:5], Y[6:4], part_p[2][6]);
part_product p0207(move_ex[2][7:6], Y[6:4], part_p[2][7]);
part_product p0208(move_ex[2][8:7], Y[6:4], part_p[2][8]);
part_product p0209(move_ex[2][9:8], Y[6:4], part_p[2][9]);
part_product p0210(move_ex[2][10:9], Y[6:4], part_p[2][10]);
part_product p0211(move_ex[2][11:10], Y[6:4], part_p[2][11]);
part_product p0212(move_ex[2][12:11], Y[6:4], part_p[2][12]);
part_product p0213(move_ex[2][13:12], Y[6:4], part_p[2][13]);
part_product p0214(move_ex[2][14:13], Y[6:4], part_p[2][14]);
part_product p0215(move_ex[2][15:14], Y[6:4], part_p[2][15]);
part_product p0216(move_ex[2][16:15], Y[6:4], part_p[2][16]);
part_product p0217(move_ex[2][17:16], Y[6:4], part_p[2][17]);
part_product p0218(move_ex[2][18:17], Y[6:4], part_p[2][18]);
part_product p0219(move_ex[2][19:18], Y[6:4], part_p[2][19]);
part_product p0220(move_ex[2][20:19], Y[6:4], part_p[2][20]);
part_product p0221(move_ex[2][21:20], Y[6:4], part_p[2][21]);
part_product p0222(move_ex[2][22:21], Y[6:4], part_p[2][22]);
part_product p0223(move_ex[2][23:22], Y[6:4], part_p[2][23]);
part_product p0224(move_ex[2][24:23], Y[6:4], part_p[2][24]);
part_product p0225(move_ex[2][25:24], Y[6:4], part_p[2][25]);
part_product p0226(move_ex[2][26:25], Y[6:4], part_p[2][26]);
part_product p0227(move_ex[2][27:26], Y[6:4], part_p[2][27]);
part_product p0228(move_ex[2][28:27], Y[6:4], part_p[2][28]);
part_product p0229(move_ex[2][29:28], Y[6:4], part_p[2][29]);
part_product p0230(move_ex[2][30:29], Y[6:4], part_p[2][30]);
part_product p0231(move_ex[2][31:30], Y[6:4], part_p[2][31]);
part_product p0232(move_ex[2][32:31], Y[6:4], part_p[2][32]);
part_product p0233(move_ex[2][33:32], Y[6:4], part_p[2][33]);
part_product p0234(move_ex[2][34:33], Y[6:4], part_p[2][34]);
part_product p0235(move_ex[2][35:34], Y[6:4], part_p[2][35]);
part_product p0236(move_ex[2][36:35], Y[6:4], part_p[2][36]);
part_product p0237(move_ex[2][37:36], Y[6:4], part_p[2][37]);
part_product p0238(move_ex[2][38:37], Y[6:4], part_p[2][38]);
part_product p0239(move_ex[2][39:38], Y[6:4], part_p[2][39]);
part_product p0240(move_ex[2][40:39], Y[6:4], part_p[2][40]);
part_product p0241(move_ex[2][41:40], Y[6:4], part_p[2][41]);
part_product p0242(move_ex[2][42:41], Y[6:4], part_p[2][42]);
part_product p0243(move_ex[2][43:42], Y[6:4], part_p[2][43]);
part_product p0244(move_ex[2][44:43], Y[6:4], part_p[2][44]);
part_product p0245(move_ex[2][45:44], Y[6:4], part_p[2][45]);
part_product p0246(move_ex[2][46:45], Y[6:4], part_p[2][46]);
part_product p0247(move_ex[2][47:46], Y[6:4], part_p[2][47]);
part_product p0248(move_ex[2][48:47], Y[6:4], part_p[2][48]);
part_product p0249(move_ex[2][49:48], Y[6:4], part_p[2][49]);
part_product p0250(move_ex[2][50:49], Y[6:4], part_p[2][50]);
part_product p0251(move_ex[2][51:50], Y[6:4], part_p[2][51]);
part_product p0252(move_ex[2][52:51], Y[6:4], part_p[2][52]);
part_product p0253(move_ex[2][53:52], Y[6:4], part_p[2][53]);
part_product p0254(move_ex[2][54:53], Y[6:4], part_p[2][54]);
part_product p0255(move_ex[2][55:54], Y[6:4], part_p[2][55]);
part_product p0256(move_ex[2][56:55], Y[6:4], part_p[2][56]);
part_product p0257(move_ex[2][57:56], Y[6:4], part_p[2][57]);
part_product p0258(move_ex[2][58:57], Y[6:4], part_p[2][58]);
part_product p0259(move_ex[2][59:58], Y[6:4], part_p[2][59]);
part_product p0260(move_ex[2][60:59], Y[6:4], part_p[2][60]);
part_product p0261(move_ex[2][61:60], Y[6:4], part_p[2][61]);
part_product p0262(move_ex[2][62:61], Y[6:4], part_p[2][62]);
part_product p0263(move_ex[2][63:62], Y[6:4], part_p[2][63]);
part_product p0264(move_ex[2][64:63], Y[6:4], part_p[2][64]);
part_product p0265(move_ex[2][65:64], Y[6:4], part_p[2][65]);
part_product p0266(move_ex[2][66:65], Y[6:4], part_p[2][66]);
part_product p0267(move_ex[2][67:66], Y[6:4], part_p[2][67]);
get_c getc2(Y[6:4], C[5:4]);

assign part_p[3][0] = 0;
assign part_p[3][1] = 0;
assign part_p[3][2] = 0;
assign part_p[3][3] = 0;
assign part_p[3][4] = 0;
assign part_p[3][5] = 0;
s_part_product sp0306(move_ex[3][6:6], Y[8:6], part_p[3][6]);
part_product p0307(move_ex[3][7:6], Y[8:6], part_p[3][7]);
part_product p0308(move_ex[3][8:7], Y[8:6], part_p[3][8]);
part_product p0309(move_ex[3][9:8], Y[8:6], part_p[3][9]);
part_product p0310(move_ex[3][10:9], Y[8:6], part_p[3][10]);
part_product p0311(move_ex[3][11:10], Y[8:6], part_p[3][11]);
part_product p0312(move_ex[3][12:11], Y[8:6], part_p[3][12]);
part_product p0313(move_ex[3][13:12], Y[8:6], part_p[3][13]);
part_product p0314(move_ex[3][14:13], Y[8:6], part_p[3][14]);
part_product p0315(move_ex[3][15:14], Y[8:6], part_p[3][15]);
part_product p0316(move_ex[3][16:15], Y[8:6], part_p[3][16]);
part_product p0317(move_ex[3][17:16], Y[8:6], part_p[3][17]);
part_product p0318(move_ex[3][18:17], Y[8:6], part_p[3][18]);
part_product p0319(move_ex[3][19:18], Y[8:6], part_p[3][19]);
part_product p0320(move_ex[3][20:19], Y[8:6], part_p[3][20]);
part_product p0321(move_ex[3][21:20], Y[8:6], part_p[3][21]);
part_product p0322(move_ex[3][22:21], Y[8:6], part_p[3][22]);
part_product p0323(move_ex[3][23:22], Y[8:6], part_p[3][23]);
part_product p0324(move_ex[3][24:23], Y[8:6], part_p[3][24]);
part_product p0325(move_ex[3][25:24], Y[8:6], part_p[3][25]);
part_product p0326(move_ex[3][26:25], Y[8:6], part_p[3][26]);
part_product p0327(move_ex[3][27:26], Y[8:6], part_p[3][27]);
part_product p0328(move_ex[3][28:27], Y[8:6], part_p[3][28]);
part_product p0329(move_ex[3][29:28], Y[8:6], part_p[3][29]);
part_product p0330(move_ex[3][30:29], Y[8:6], part_p[3][30]);
part_product p0331(move_ex[3][31:30], Y[8:6], part_p[3][31]);
part_product p0332(move_ex[3][32:31], Y[8:6], part_p[3][32]);
part_product p0333(move_ex[3][33:32], Y[8:6], part_p[3][33]);
part_product p0334(move_ex[3][34:33], Y[8:6], part_p[3][34]);
part_product p0335(move_ex[3][35:34], Y[8:6], part_p[3][35]);
part_product p0336(move_ex[3][36:35], Y[8:6], part_p[3][36]);
part_product p0337(move_ex[3][37:36], Y[8:6], part_p[3][37]);
part_product p0338(move_ex[3][38:37], Y[8:6], part_p[3][38]);
part_product p0339(move_ex[3][39:38], Y[8:6], part_p[3][39]);
part_product p0340(move_ex[3][40:39], Y[8:6], part_p[3][40]);
part_product p0341(move_ex[3][41:40], Y[8:6], part_p[3][41]);
part_product p0342(move_ex[3][42:41], Y[8:6], part_p[3][42]);
part_product p0343(move_ex[3][43:42], Y[8:6], part_p[3][43]);
part_product p0344(move_ex[3][44:43], Y[8:6], part_p[3][44]);
part_product p0345(move_ex[3][45:44], Y[8:6], part_p[3][45]);
part_product p0346(move_ex[3][46:45], Y[8:6], part_p[3][46]);
part_product p0347(move_ex[3][47:46], Y[8:6], part_p[3][47]);
part_product p0348(move_ex[3][48:47], Y[8:6], part_p[3][48]);
part_product p0349(move_ex[3][49:48], Y[8:6], part_p[3][49]);
part_product p0350(move_ex[3][50:49], Y[8:6], part_p[3][50]);
part_product p0351(move_ex[3][51:50], Y[8:6], part_p[3][51]);
part_product p0352(move_ex[3][52:51], Y[8:6], part_p[3][52]);
part_product p0353(move_ex[3][53:52], Y[8:6], part_p[3][53]);
part_product p0354(move_ex[3][54:53], Y[8:6], part_p[3][54]);
part_product p0355(move_ex[3][55:54], Y[8:6], part_p[3][55]);
part_product p0356(move_ex[3][56:55], Y[8:6], part_p[3][56]);
part_product p0357(move_ex[3][57:56], Y[8:6], part_p[3][57]);
part_product p0358(move_ex[3][58:57], Y[8:6], part_p[3][58]);
part_product p0359(move_ex[3][59:58], Y[8:6], part_p[3][59]);
part_product p0360(move_ex[3][60:59], Y[8:6], part_p[3][60]);
part_product p0361(move_ex[3][61:60], Y[8:6], part_p[3][61]);
part_product p0362(move_ex[3][62:61], Y[8:6], part_p[3][62]);
part_product p0363(move_ex[3][63:62], Y[8:6], part_p[3][63]);
part_product p0364(move_ex[3][64:63], Y[8:6], part_p[3][64]);
part_product p0365(move_ex[3][65:64], Y[8:6], part_p[3][65]);
part_product p0366(move_ex[3][66:65], Y[8:6], part_p[3][66]);
part_product p0367(move_ex[3][67:66], Y[8:6], part_p[3][67]);
get_c getc3(Y[8:6], C[7:6]);

assign part_p[4][0] = 0;
assign part_p[4][1] = 0;
assign part_p[4][2] = 0;
assign part_p[4][3] = 0;
assign part_p[4][4] = 0;
assign part_p[4][5] = 0;
assign part_p[4][6] = 0;
assign part_p[4][7] = 0;
s_part_product sp0408(move_ex[4][8:8], Y[10:8], part_p[4][8]);
part_product p0409(move_ex[4][9:8], Y[10:8], part_p[4][9]);
part_product p0410(move_ex[4][10:9], Y[10:8], part_p[4][10]);
part_product p0411(move_ex[4][11:10], Y[10:8], part_p[4][11]);
part_product p0412(move_ex[4][12:11], Y[10:8], part_p[4][12]);
part_product p0413(move_ex[4][13:12], Y[10:8], part_p[4][13]);
part_product p0414(move_ex[4][14:13], Y[10:8], part_p[4][14]);
part_product p0415(move_ex[4][15:14], Y[10:8], part_p[4][15]);
part_product p0416(move_ex[4][16:15], Y[10:8], part_p[4][16]);
part_product p0417(move_ex[4][17:16], Y[10:8], part_p[4][17]);
part_product p0418(move_ex[4][18:17], Y[10:8], part_p[4][18]);
part_product p0419(move_ex[4][19:18], Y[10:8], part_p[4][19]);
part_product p0420(move_ex[4][20:19], Y[10:8], part_p[4][20]);
part_product p0421(move_ex[4][21:20], Y[10:8], part_p[4][21]);
part_product p0422(move_ex[4][22:21], Y[10:8], part_p[4][22]);
part_product p0423(move_ex[4][23:22], Y[10:8], part_p[4][23]);
part_product p0424(move_ex[4][24:23], Y[10:8], part_p[4][24]);
part_product p0425(move_ex[4][25:24], Y[10:8], part_p[4][25]);
part_product p0426(move_ex[4][26:25], Y[10:8], part_p[4][26]);
part_product p0427(move_ex[4][27:26], Y[10:8], part_p[4][27]);
part_product p0428(move_ex[4][28:27], Y[10:8], part_p[4][28]);
part_product p0429(move_ex[4][29:28], Y[10:8], part_p[4][29]);
part_product p0430(move_ex[4][30:29], Y[10:8], part_p[4][30]);
part_product p0431(move_ex[4][31:30], Y[10:8], part_p[4][31]);
part_product p0432(move_ex[4][32:31], Y[10:8], part_p[4][32]);
part_product p0433(move_ex[4][33:32], Y[10:8], part_p[4][33]);
part_product p0434(move_ex[4][34:33], Y[10:8], part_p[4][34]);
part_product p0435(move_ex[4][35:34], Y[10:8], part_p[4][35]);
part_product p0436(move_ex[4][36:35], Y[10:8], part_p[4][36]);
part_product p0437(move_ex[4][37:36], Y[10:8], part_p[4][37]);
part_product p0438(move_ex[4][38:37], Y[10:8], part_p[4][38]);
part_product p0439(move_ex[4][39:38], Y[10:8], part_p[4][39]);
part_product p0440(move_ex[4][40:39], Y[10:8], part_p[4][40]);
part_product p0441(move_ex[4][41:40], Y[10:8], part_p[4][41]);
part_product p0442(move_ex[4][42:41], Y[10:8], part_p[4][42]);
part_product p0443(move_ex[4][43:42], Y[10:8], part_p[4][43]);
part_product p0444(move_ex[4][44:43], Y[10:8], part_p[4][44]);
part_product p0445(move_ex[4][45:44], Y[10:8], part_p[4][45]);
part_product p0446(move_ex[4][46:45], Y[10:8], part_p[4][46]);
part_product p0447(move_ex[4][47:46], Y[10:8], part_p[4][47]);
part_product p0448(move_ex[4][48:47], Y[10:8], part_p[4][48]);
part_product p0449(move_ex[4][49:48], Y[10:8], part_p[4][49]);
part_product p0450(move_ex[4][50:49], Y[10:8], part_p[4][50]);
part_product p0451(move_ex[4][51:50], Y[10:8], part_p[4][51]);
part_product p0452(move_ex[4][52:51], Y[10:8], part_p[4][52]);
part_product p0453(move_ex[4][53:52], Y[10:8], part_p[4][53]);
part_product p0454(move_ex[4][54:53], Y[10:8], part_p[4][54]);
part_product p0455(move_ex[4][55:54], Y[10:8], part_p[4][55]);
part_product p0456(move_ex[4][56:55], Y[10:8], part_p[4][56]);
part_product p0457(move_ex[4][57:56], Y[10:8], part_p[4][57]);
part_product p0458(move_ex[4][58:57], Y[10:8], part_p[4][58]);
part_product p0459(move_ex[4][59:58], Y[10:8], part_p[4][59]);
part_product p0460(move_ex[4][60:59], Y[10:8], part_p[4][60]);
part_product p0461(move_ex[4][61:60], Y[10:8], part_p[4][61]);
part_product p0462(move_ex[4][62:61], Y[10:8], part_p[4][62]);
part_product p0463(move_ex[4][63:62], Y[10:8], part_p[4][63]);
part_product p0464(move_ex[4][64:63], Y[10:8], part_p[4][64]);
part_product p0465(move_ex[4][65:64], Y[10:8], part_p[4][65]);
part_product p0466(move_ex[4][66:65], Y[10:8], part_p[4][66]);
part_product p0467(move_ex[4][67:66], Y[10:8], part_p[4][67]);
get_c getc4(Y[10:8], C[9:8]);

assign part_p[5][0] = 0;
assign part_p[5][1] = 0;
assign part_p[5][2] = 0;
assign part_p[5][3] = 0;
assign part_p[5][4] = 0;
assign part_p[5][5] = 0;
assign part_p[5][6] = 0;
assign part_p[5][7] = 0;
assign part_p[5][8] = 0;
assign part_p[5][9] = 0;
s_part_product sp0510(move_ex[5][10:10], Y[12:10], part_p[5][10]);
part_product p0511(move_ex[5][11:10], Y[12:10], part_p[5][11]);
part_product p0512(move_ex[5][12:11], Y[12:10], part_p[5][12]);
part_product p0513(move_ex[5][13:12], Y[12:10], part_p[5][13]);
part_product p0514(move_ex[5][14:13], Y[12:10], part_p[5][14]);
part_product p0515(move_ex[5][15:14], Y[12:10], part_p[5][15]);
part_product p0516(move_ex[5][16:15], Y[12:10], part_p[5][16]);
part_product p0517(move_ex[5][17:16], Y[12:10], part_p[5][17]);
part_product p0518(move_ex[5][18:17], Y[12:10], part_p[5][18]);
part_product p0519(move_ex[5][19:18], Y[12:10], part_p[5][19]);
part_product p0520(move_ex[5][20:19], Y[12:10], part_p[5][20]);
part_product p0521(move_ex[5][21:20], Y[12:10], part_p[5][21]);
part_product p0522(move_ex[5][22:21], Y[12:10], part_p[5][22]);
part_product p0523(move_ex[5][23:22], Y[12:10], part_p[5][23]);
part_product p0524(move_ex[5][24:23], Y[12:10], part_p[5][24]);
part_product p0525(move_ex[5][25:24], Y[12:10], part_p[5][25]);
part_product p0526(move_ex[5][26:25], Y[12:10], part_p[5][26]);
part_product p0527(move_ex[5][27:26], Y[12:10], part_p[5][27]);
part_product p0528(move_ex[5][28:27], Y[12:10], part_p[5][28]);
part_product p0529(move_ex[5][29:28], Y[12:10], part_p[5][29]);
part_product p0530(move_ex[5][30:29], Y[12:10], part_p[5][30]);
part_product p0531(move_ex[5][31:30], Y[12:10], part_p[5][31]);
part_product p0532(move_ex[5][32:31], Y[12:10], part_p[5][32]);
part_product p0533(move_ex[5][33:32], Y[12:10], part_p[5][33]);
part_product p0534(move_ex[5][34:33], Y[12:10], part_p[5][34]);
part_product p0535(move_ex[5][35:34], Y[12:10], part_p[5][35]);
part_product p0536(move_ex[5][36:35], Y[12:10], part_p[5][36]);
part_product p0537(move_ex[5][37:36], Y[12:10], part_p[5][37]);
part_product p0538(move_ex[5][38:37], Y[12:10], part_p[5][38]);
part_product p0539(move_ex[5][39:38], Y[12:10], part_p[5][39]);
part_product p0540(move_ex[5][40:39], Y[12:10], part_p[5][40]);
part_product p0541(move_ex[5][41:40], Y[12:10], part_p[5][41]);
part_product p0542(move_ex[5][42:41], Y[12:10], part_p[5][42]);
part_product p0543(move_ex[5][43:42], Y[12:10], part_p[5][43]);
part_product p0544(move_ex[5][44:43], Y[12:10], part_p[5][44]);
part_product p0545(move_ex[5][45:44], Y[12:10], part_p[5][45]);
part_product p0546(move_ex[5][46:45], Y[12:10], part_p[5][46]);
part_product p0547(move_ex[5][47:46], Y[12:10], part_p[5][47]);
part_product p0548(move_ex[5][48:47], Y[12:10], part_p[5][48]);
part_product p0549(move_ex[5][49:48], Y[12:10], part_p[5][49]);
part_product p0550(move_ex[5][50:49], Y[12:10], part_p[5][50]);
part_product p0551(move_ex[5][51:50], Y[12:10], part_p[5][51]);
part_product p0552(move_ex[5][52:51], Y[12:10], part_p[5][52]);
part_product p0553(move_ex[5][53:52], Y[12:10], part_p[5][53]);
part_product p0554(move_ex[5][54:53], Y[12:10], part_p[5][54]);
part_product p0555(move_ex[5][55:54], Y[12:10], part_p[5][55]);
part_product p0556(move_ex[5][56:55], Y[12:10], part_p[5][56]);
part_product p0557(move_ex[5][57:56], Y[12:10], part_p[5][57]);
part_product p0558(move_ex[5][58:57], Y[12:10], part_p[5][58]);
part_product p0559(move_ex[5][59:58], Y[12:10], part_p[5][59]);
part_product p0560(move_ex[5][60:59], Y[12:10], part_p[5][60]);
part_product p0561(move_ex[5][61:60], Y[12:10], part_p[5][61]);
part_product p0562(move_ex[5][62:61], Y[12:10], part_p[5][62]);
part_product p0563(move_ex[5][63:62], Y[12:10], part_p[5][63]);
part_product p0564(move_ex[5][64:63], Y[12:10], part_p[5][64]);
part_product p0565(move_ex[5][65:64], Y[12:10], part_p[5][65]);
part_product p0566(move_ex[5][66:65], Y[12:10], part_p[5][66]);
part_product p0567(move_ex[5][67:66], Y[12:10], part_p[5][67]);
get_c getc5(Y[12:10], C[11:10]);

assign part_p[6][0] = 0;
assign part_p[6][1] = 0;
assign part_p[6][2] = 0;
assign part_p[6][3] = 0;
assign part_p[6][4] = 0;
assign part_p[6][5] = 0;
assign part_p[6][6] = 0;
assign part_p[6][7] = 0;
assign part_p[6][8] = 0;
assign part_p[6][9] = 0;
assign part_p[6][10] = 0;
assign part_p[6][11] = 0;
s_part_product sp0612(move_ex[6][12:12], Y[14:12], part_p[6][12]);
part_product p0613(move_ex[6][13:12], Y[14:12], part_p[6][13]);
part_product p0614(move_ex[6][14:13], Y[14:12], part_p[6][14]);
part_product p0615(move_ex[6][15:14], Y[14:12], part_p[6][15]);
part_product p0616(move_ex[6][16:15], Y[14:12], part_p[6][16]);
part_product p0617(move_ex[6][17:16], Y[14:12], part_p[6][17]);
part_product p0618(move_ex[6][18:17], Y[14:12], part_p[6][18]);
part_product p0619(move_ex[6][19:18], Y[14:12], part_p[6][19]);
part_product p0620(move_ex[6][20:19], Y[14:12], part_p[6][20]);
part_product p0621(move_ex[6][21:20], Y[14:12], part_p[6][21]);
part_product p0622(move_ex[6][22:21], Y[14:12], part_p[6][22]);
part_product p0623(move_ex[6][23:22], Y[14:12], part_p[6][23]);
part_product p0624(move_ex[6][24:23], Y[14:12], part_p[6][24]);
part_product p0625(move_ex[6][25:24], Y[14:12], part_p[6][25]);
part_product p0626(move_ex[6][26:25], Y[14:12], part_p[6][26]);
part_product p0627(move_ex[6][27:26], Y[14:12], part_p[6][27]);
part_product p0628(move_ex[6][28:27], Y[14:12], part_p[6][28]);
part_product p0629(move_ex[6][29:28], Y[14:12], part_p[6][29]);
part_product p0630(move_ex[6][30:29], Y[14:12], part_p[6][30]);
part_product p0631(move_ex[6][31:30], Y[14:12], part_p[6][31]);
part_product p0632(move_ex[6][32:31], Y[14:12], part_p[6][32]);
part_product p0633(move_ex[6][33:32], Y[14:12], part_p[6][33]);
part_product p0634(move_ex[6][34:33], Y[14:12], part_p[6][34]);
part_product p0635(move_ex[6][35:34], Y[14:12], part_p[6][35]);
part_product p0636(move_ex[6][36:35], Y[14:12], part_p[6][36]);
part_product p0637(move_ex[6][37:36], Y[14:12], part_p[6][37]);
part_product p0638(move_ex[6][38:37], Y[14:12], part_p[6][38]);
part_product p0639(move_ex[6][39:38], Y[14:12], part_p[6][39]);
part_product p0640(move_ex[6][40:39], Y[14:12], part_p[6][40]);
part_product p0641(move_ex[6][41:40], Y[14:12], part_p[6][41]);
part_product p0642(move_ex[6][42:41], Y[14:12], part_p[6][42]);
part_product p0643(move_ex[6][43:42], Y[14:12], part_p[6][43]);
part_product p0644(move_ex[6][44:43], Y[14:12], part_p[6][44]);
part_product p0645(move_ex[6][45:44], Y[14:12], part_p[6][45]);
part_product p0646(move_ex[6][46:45], Y[14:12], part_p[6][46]);
part_product p0647(move_ex[6][47:46], Y[14:12], part_p[6][47]);
part_product p0648(move_ex[6][48:47], Y[14:12], part_p[6][48]);
part_product p0649(move_ex[6][49:48], Y[14:12], part_p[6][49]);
part_product p0650(move_ex[6][50:49], Y[14:12], part_p[6][50]);
part_product p0651(move_ex[6][51:50], Y[14:12], part_p[6][51]);
part_product p0652(move_ex[6][52:51], Y[14:12], part_p[6][52]);
part_product p0653(move_ex[6][53:52], Y[14:12], part_p[6][53]);
part_product p0654(move_ex[6][54:53], Y[14:12], part_p[6][54]);
part_product p0655(move_ex[6][55:54], Y[14:12], part_p[6][55]);
part_product p0656(move_ex[6][56:55], Y[14:12], part_p[6][56]);
part_product p0657(move_ex[6][57:56], Y[14:12], part_p[6][57]);
part_product p0658(move_ex[6][58:57], Y[14:12], part_p[6][58]);
part_product p0659(move_ex[6][59:58], Y[14:12], part_p[6][59]);
part_product p0660(move_ex[6][60:59], Y[14:12], part_p[6][60]);
part_product p0661(move_ex[6][61:60], Y[14:12], part_p[6][61]);
part_product p0662(move_ex[6][62:61], Y[14:12], part_p[6][62]);
part_product p0663(move_ex[6][63:62], Y[14:12], part_p[6][63]);
part_product p0664(move_ex[6][64:63], Y[14:12], part_p[6][64]);
part_product p0665(move_ex[6][65:64], Y[14:12], part_p[6][65]);
part_product p0666(move_ex[6][66:65], Y[14:12], part_p[6][66]);
part_product p0667(move_ex[6][67:66], Y[14:12], part_p[6][67]);
get_c getc6(Y[14:12], C[13:12]);

assign part_p[7][0] = 0;
assign part_p[7][1] = 0;
assign part_p[7][2] = 0;
assign part_p[7][3] = 0;
assign part_p[7][4] = 0;
assign part_p[7][5] = 0;
assign part_p[7][6] = 0;
assign part_p[7][7] = 0;
assign part_p[7][8] = 0;
assign part_p[7][9] = 0;
assign part_p[7][10] = 0;
assign part_p[7][11] = 0;
assign part_p[7][12] = 0;
assign part_p[7][13] = 0;
s_part_product sp0714(move_ex[7][14:14], Y[16:14], part_p[7][14]);
part_product p0715(move_ex[7][15:14], Y[16:14], part_p[7][15]);
part_product p0716(move_ex[7][16:15], Y[16:14], part_p[7][16]);
part_product p0717(move_ex[7][17:16], Y[16:14], part_p[7][17]);
part_product p0718(move_ex[7][18:17], Y[16:14], part_p[7][18]);
part_product p0719(move_ex[7][19:18], Y[16:14], part_p[7][19]);
part_product p0720(move_ex[7][20:19], Y[16:14], part_p[7][20]);
part_product p0721(move_ex[7][21:20], Y[16:14], part_p[7][21]);
part_product p0722(move_ex[7][22:21], Y[16:14], part_p[7][22]);
part_product p0723(move_ex[7][23:22], Y[16:14], part_p[7][23]);
part_product p0724(move_ex[7][24:23], Y[16:14], part_p[7][24]);
part_product p0725(move_ex[7][25:24], Y[16:14], part_p[7][25]);
part_product p0726(move_ex[7][26:25], Y[16:14], part_p[7][26]);
part_product p0727(move_ex[7][27:26], Y[16:14], part_p[7][27]);
part_product p0728(move_ex[7][28:27], Y[16:14], part_p[7][28]);
part_product p0729(move_ex[7][29:28], Y[16:14], part_p[7][29]);
part_product p0730(move_ex[7][30:29], Y[16:14], part_p[7][30]);
part_product p0731(move_ex[7][31:30], Y[16:14], part_p[7][31]);
part_product p0732(move_ex[7][32:31], Y[16:14], part_p[7][32]);
part_product p0733(move_ex[7][33:32], Y[16:14], part_p[7][33]);
part_product p0734(move_ex[7][34:33], Y[16:14], part_p[7][34]);
part_product p0735(move_ex[7][35:34], Y[16:14], part_p[7][35]);
part_product p0736(move_ex[7][36:35], Y[16:14], part_p[7][36]);
part_product p0737(move_ex[7][37:36], Y[16:14], part_p[7][37]);
part_product p0738(move_ex[7][38:37], Y[16:14], part_p[7][38]);
part_product p0739(move_ex[7][39:38], Y[16:14], part_p[7][39]);
part_product p0740(move_ex[7][40:39], Y[16:14], part_p[7][40]);
part_product p0741(move_ex[7][41:40], Y[16:14], part_p[7][41]);
part_product p0742(move_ex[7][42:41], Y[16:14], part_p[7][42]);
part_product p0743(move_ex[7][43:42], Y[16:14], part_p[7][43]);
part_product p0744(move_ex[7][44:43], Y[16:14], part_p[7][44]);
part_product p0745(move_ex[7][45:44], Y[16:14], part_p[7][45]);
part_product p0746(move_ex[7][46:45], Y[16:14], part_p[7][46]);
part_product p0747(move_ex[7][47:46], Y[16:14], part_p[7][47]);
part_product p0748(move_ex[7][48:47], Y[16:14], part_p[7][48]);
part_product p0749(move_ex[7][49:48], Y[16:14], part_p[7][49]);
part_product p0750(move_ex[7][50:49], Y[16:14], part_p[7][50]);
part_product p0751(move_ex[7][51:50], Y[16:14], part_p[7][51]);
part_product p0752(move_ex[7][52:51], Y[16:14], part_p[7][52]);
part_product p0753(move_ex[7][53:52], Y[16:14], part_p[7][53]);
part_product p0754(move_ex[7][54:53], Y[16:14], part_p[7][54]);
part_product p0755(move_ex[7][55:54], Y[16:14], part_p[7][55]);
part_product p0756(move_ex[7][56:55], Y[16:14], part_p[7][56]);
part_product p0757(move_ex[7][57:56], Y[16:14], part_p[7][57]);
part_product p0758(move_ex[7][58:57], Y[16:14], part_p[7][58]);
part_product p0759(move_ex[7][59:58], Y[16:14], part_p[7][59]);
part_product p0760(move_ex[7][60:59], Y[16:14], part_p[7][60]);
part_product p0761(move_ex[7][61:60], Y[16:14], part_p[7][61]);
part_product p0762(move_ex[7][62:61], Y[16:14], part_p[7][62]);
part_product p0763(move_ex[7][63:62], Y[16:14], part_p[7][63]);
part_product p0764(move_ex[7][64:63], Y[16:14], part_p[7][64]);
part_product p0765(move_ex[7][65:64], Y[16:14], part_p[7][65]);
part_product p0766(move_ex[7][66:65], Y[16:14], part_p[7][66]);
part_product p0767(move_ex[7][67:66], Y[16:14], part_p[7][67]);
get_c getc7(Y[16:14], C[15:14]);

assign part_p[8][0] = 0;
assign part_p[8][1] = 0;
assign part_p[8][2] = 0;
assign part_p[8][3] = 0;
assign part_p[8][4] = 0;
assign part_p[8][5] = 0;
assign part_p[8][6] = 0;
assign part_p[8][7] = 0;
assign part_p[8][8] = 0;
assign part_p[8][9] = 0;
assign part_p[8][10] = 0;
assign part_p[8][11] = 0;
assign part_p[8][12] = 0;
assign part_p[8][13] = 0;
assign part_p[8][14] = 0;
assign part_p[8][15] = 0;
s_part_product sp0816(move_ex[8][16:16], Y[18:16], part_p[8][16]);
part_product p0817(move_ex[8][17:16], Y[18:16], part_p[8][17]);
part_product p0818(move_ex[8][18:17], Y[18:16], part_p[8][18]);
part_product p0819(move_ex[8][19:18], Y[18:16], part_p[8][19]);
part_product p0820(move_ex[8][20:19], Y[18:16], part_p[8][20]);
part_product p0821(move_ex[8][21:20], Y[18:16], part_p[8][21]);
part_product p0822(move_ex[8][22:21], Y[18:16], part_p[8][22]);
part_product p0823(move_ex[8][23:22], Y[18:16], part_p[8][23]);
part_product p0824(move_ex[8][24:23], Y[18:16], part_p[8][24]);
part_product p0825(move_ex[8][25:24], Y[18:16], part_p[8][25]);
part_product p0826(move_ex[8][26:25], Y[18:16], part_p[8][26]);
part_product p0827(move_ex[8][27:26], Y[18:16], part_p[8][27]);
part_product p0828(move_ex[8][28:27], Y[18:16], part_p[8][28]);
part_product p0829(move_ex[8][29:28], Y[18:16], part_p[8][29]);
part_product p0830(move_ex[8][30:29], Y[18:16], part_p[8][30]);
part_product p0831(move_ex[8][31:30], Y[18:16], part_p[8][31]);
part_product p0832(move_ex[8][32:31], Y[18:16], part_p[8][32]);
part_product p0833(move_ex[8][33:32], Y[18:16], part_p[8][33]);
part_product p0834(move_ex[8][34:33], Y[18:16], part_p[8][34]);
part_product p0835(move_ex[8][35:34], Y[18:16], part_p[8][35]);
part_product p0836(move_ex[8][36:35], Y[18:16], part_p[8][36]);
part_product p0837(move_ex[8][37:36], Y[18:16], part_p[8][37]);
part_product p0838(move_ex[8][38:37], Y[18:16], part_p[8][38]);
part_product p0839(move_ex[8][39:38], Y[18:16], part_p[8][39]);
part_product p0840(move_ex[8][40:39], Y[18:16], part_p[8][40]);
part_product p0841(move_ex[8][41:40], Y[18:16], part_p[8][41]);
part_product p0842(move_ex[8][42:41], Y[18:16], part_p[8][42]);
part_product p0843(move_ex[8][43:42], Y[18:16], part_p[8][43]);
part_product p0844(move_ex[8][44:43], Y[18:16], part_p[8][44]);
part_product p0845(move_ex[8][45:44], Y[18:16], part_p[8][45]);
part_product p0846(move_ex[8][46:45], Y[18:16], part_p[8][46]);
part_product p0847(move_ex[8][47:46], Y[18:16], part_p[8][47]);
part_product p0848(move_ex[8][48:47], Y[18:16], part_p[8][48]);
part_product p0849(move_ex[8][49:48], Y[18:16], part_p[8][49]);
part_product p0850(move_ex[8][50:49], Y[18:16], part_p[8][50]);
part_product p0851(move_ex[8][51:50], Y[18:16], part_p[8][51]);
part_product p0852(move_ex[8][52:51], Y[18:16], part_p[8][52]);
part_product p0853(move_ex[8][53:52], Y[18:16], part_p[8][53]);
part_product p0854(move_ex[8][54:53], Y[18:16], part_p[8][54]);
part_product p0855(move_ex[8][55:54], Y[18:16], part_p[8][55]);
part_product p0856(move_ex[8][56:55], Y[18:16], part_p[8][56]);
part_product p0857(move_ex[8][57:56], Y[18:16], part_p[8][57]);
part_product p0858(move_ex[8][58:57], Y[18:16], part_p[8][58]);
part_product p0859(move_ex[8][59:58], Y[18:16], part_p[8][59]);
part_product p0860(move_ex[8][60:59], Y[18:16], part_p[8][60]);
part_product p0861(move_ex[8][61:60], Y[18:16], part_p[8][61]);
part_product p0862(move_ex[8][62:61], Y[18:16], part_p[8][62]);
part_product p0863(move_ex[8][63:62], Y[18:16], part_p[8][63]);
part_product p0864(move_ex[8][64:63], Y[18:16], part_p[8][64]);
part_product p0865(move_ex[8][65:64], Y[18:16], part_p[8][65]);
part_product p0866(move_ex[8][66:65], Y[18:16], part_p[8][66]);
part_product p0867(move_ex[8][67:66], Y[18:16], part_p[8][67]);
get_c getc8(Y[18:16], C[17:16]);

assign part_p[9][0] = 0;
assign part_p[9][1] = 0;
assign part_p[9][2] = 0;
assign part_p[9][3] = 0;
assign part_p[9][4] = 0;
assign part_p[9][5] = 0;
assign part_p[9][6] = 0;
assign part_p[9][7] = 0;
assign part_p[9][8] = 0;
assign part_p[9][9] = 0;
assign part_p[9][10] = 0;
assign part_p[9][11] = 0;
assign part_p[9][12] = 0;
assign part_p[9][13] = 0;
assign part_p[9][14] = 0;
assign part_p[9][15] = 0;
assign part_p[9][16] = 0;
assign part_p[9][17] = 0;
s_part_product sp0918(move_ex[9][18:18], Y[20:18], part_p[9][18]);
part_product p0919(move_ex[9][19:18], Y[20:18], part_p[9][19]);
part_product p0920(move_ex[9][20:19], Y[20:18], part_p[9][20]);
part_product p0921(move_ex[9][21:20], Y[20:18], part_p[9][21]);
part_product p0922(move_ex[9][22:21], Y[20:18], part_p[9][22]);
part_product p0923(move_ex[9][23:22], Y[20:18], part_p[9][23]);
part_product p0924(move_ex[9][24:23], Y[20:18], part_p[9][24]);
part_product p0925(move_ex[9][25:24], Y[20:18], part_p[9][25]);
part_product p0926(move_ex[9][26:25], Y[20:18], part_p[9][26]);
part_product p0927(move_ex[9][27:26], Y[20:18], part_p[9][27]);
part_product p0928(move_ex[9][28:27], Y[20:18], part_p[9][28]);
part_product p0929(move_ex[9][29:28], Y[20:18], part_p[9][29]);
part_product p0930(move_ex[9][30:29], Y[20:18], part_p[9][30]);
part_product p0931(move_ex[9][31:30], Y[20:18], part_p[9][31]);
part_product p0932(move_ex[9][32:31], Y[20:18], part_p[9][32]);
part_product p0933(move_ex[9][33:32], Y[20:18], part_p[9][33]);
part_product p0934(move_ex[9][34:33], Y[20:18], part_p[9][34]);
part_product p0935(move_ex[9][35:34], Y[20:18], part_p[9][35]);
part_product p0936(move_ex[9][36:35], Y[20:18], part_p[9][36]);
part_product p0937(move_ex[9][37:36], Y[20:18], part_p[9][37]);
part_product p0938(move_ex[9][38:37], Y[20:18], part_p[9][38]);
part_product p0939(move_ex[9][39:38], Y[20:18], part_p[9][39]);
part_product p0940(move_ex[9][40:39], Y[20:18], part_p[9][40]);
part_product p0941(move_ex[9][41:40], Y[20:18], part_p[9][41]);
part_product p0942(move_ex[9][42:41], Y[20:18], part_p[9][42]);
part_product p0943(move_ex[9][43:42], Y[20:18], part_p[9][43]);
part_product p0944(move_ex[9][44:43], Y[20:18], part_p[9][44]);
part_product p0945(move_ex[9][45:44], Y[20:18], part_p[9][45]);
part_product p0946(move_ex[9][46:45], Y[20:18], part_p[9][46]);
part_product p0947(move_ex[9][47:46], Y[20:18], part_p[9][47]);
part_product p0948(move_ex[9][48:47], Y[20:18], part_p[9][48]);
part_product p0949(move_ex[9][49:48], Y[20:18], part_p[9][49]);
part_product p0950(move_ex[9][50:49], Y[20:18], part_p[9][50]);
part_product p0951(move_ex[9][51:50], Y[20:18], part_p[9][51]);
part_product p0952(move_ex[9][52:51], Y[20:18], part_p[9][52]);
part_product p0953(move_ex[9][53:52], Y[20:18], part_p[9][53]);
part_product p0954(move_ex[9][54:53], Y[20:18], part_p[9][54]);
part_product p0955(move_ex[9][55:54], Y[20:18], part_p[9][55]);
part_product p0956(move_ex[9][56:55], Y[20:18], part_p[9][56]);
part_product p0957(move_ex[9][57:56], Y[20:18], part_p[9][57]);
part_product p0958(move_ex[9][58:57], Y[20:18], part_p[9][58]);
part_product p0959(move_ex[9][59:58], Y[20:18], part_p[9][59]);
part_product p0960(move_ex[9][60:59], Y[20:18], part_p[9][60]);
part_product p0961(move_ex[9][61:60], Y[20:18], part_p[9][61]);
part_product p0962(move_ex[9][62:61], Y[20:18], part_p[9][62]);
part_product p0963(move_ex[9][63:62], Y[20:18], part_p[9][63]);
part_product p0964(move_ex[9][64:63], Y[20:18], part_p[9][64]);
part_product p0965(move_ex[9][65:64], Y[20:18], part_p[9][65]);
part_product p0966(move_ex[9][66:65], Y[20:18], part_p[9][66]);
part_product p0967(move_ex[9][67:66], Y[20:18], part_p[9][67]);
get_c getc9(Y[20:18], C[19:18]);

assign part_p[10][0] = 0;
assign part_p[10][1] = 0;
assign part_p[10][2] = 0;
assign part_p[10][3] = 0;
assign part_p[10][4] = 0;
assign part_p[10][5] = 0;
assign part_p[10][6] = 0;
assign part_p[10][7] = 0;
assign part_p[10][8] = 0;
assign part_p[10][9] = 0;
assign part_p[10][10] = 0;
assign part_p[10][11] = 0;
assign part_p[10][12] = 0;
assign part_p[10][13] = 0;
assign part_p[10][14] = 0;
assign part_p[10][15] = 0;
assign part_p[10][16] = 0;
assign part_p[10][17] = 0;
assign part_p[10][18] = 0;
assign part_p[10][19] = 0;
s_part_product sp1020(move_ex[10][20:20], Y[22:20], part_p[10][20]);
part_product p1021(move_ex[10][21:20], Y[22:20], part_p[10][21]);
part_product p1022(move_ex[10][22:21], Y[22:20], part_p[10][22]);
part_product p1023(move_ex[10][23:22], Y[22:20], part_p[10][23]);
part_product p1024(move_ex[10][24:23], Y[22:20], part_p[10][24]);
part_product p1025(move_ex[10][25:24], Y[22:20], part_p[10][25]);
part_product p1026(move_ex[10][26:25], Y[22:20], part_p[10][26]);
part_product p1027(move_ex[10][27:26], Y[22:20], part_p[10][27]);
part_product p1028(move_ex[10][28:27], Y[22:20], part_p[10][28]);
part_product p1029(move_ex[10][29:28], Y[22:20], part_p[10][29]);
part_product p1030(move_ex[10][30:29], Y[22:20], part_p[10][30]);
part_product p1031(move_ex[10][31:30], Y[22:20], part_p[10][31]);
part_product p1032(move_ex[10][32:31], Y[22:20], part_p[10][32]);
part_product p1033(move_ex[10][33:32], Y[22:20], part_p[10][33]);
part_product p1034(move_ex[10][34:33], Y[22:20], part_p[10][34]);
part_product p1035(move_ex[10][35:34], Y[22:20], part_p[10][35]);
part_product p1036(move_ex[10][36:35], Y[22:20], part_p[10][36]);
part_product p1037(move_ex[10][37:36], Y[22:20], part_p[10][37]);
part_product p1038(move_ex[10][38:37], Y[22:20], part_p[10][38]);
part_product p1039(move_ex[10][39:38], Y[22:20], part_p[10][39]);
part_product p1040(move_ex[10][40:39], Y[22:20], part_p[10][40]);
part_product p1041(move_ex[10][41:40], Y[22:20], part_p[10][41]);
part_product p1042(move_ex[10][42:41], Y[22:20], part_p[10][42]);
part_product p1043(move_ex[10][43:42], Y[22:20], part_p[10][43]);
part_product p1044(move_ex[10][44:43], Y[22:20], part_p[10][44]);
part_product p1045(move_ex[10][45:44], Y[22:20], part_p[10][45]);
part_product p1046(move_ex[10][46:45], Y[22:20], part_p[10][46]);
part_product p1047(move_ex[10][47:46], Y[22:20], part_p[10][47]);
part_product p1048(move_ex[10][48:47], Y[22:20], part_p[10][48]);
part_product p1049(move_ex[10][49:48], Y[22:20], part_p[10][49]);
part_product p1050(move_ex[10][50:49], Y[22:20], part_p[10][50]);
part_product p1051(move_ex[10][51:50], Y[22:20], part_p[10][51]);
part_product p1052(move_ex[10][52:51], Y[22:20], part_p[10][52]);
part_product p1053(move_ex[10][53:52], Y[22:20], part_p[10][53]);
part_product p1054(move_ex[10][54:53], Y[22:20], part_p[10][54]);
part_product p1055(move_ex[10][55:54], Y[22:20], part_p[10][55]);
part_product p1056(move_ex[10][56:55], Y[22:20], part_p[10][56]);
part_product p1057(move_ex[10][57:56], Y[22:20], part_p[10][57]);
part_product p1058(move_ex[10][58:57], Y[22:20], part_p[10][58]);
part_product p1059(move_ex[10][59:58], Y[22:20], part_p[10][59]);
part_product p1060(move_ex[10][60:59], Y[22:20], part_p[10][60]);
part_product p1061(move_ex[10][61:60], Y[22:20], part_p[10][61]);
part_product p1062(move_ex[10][62:61], Y[22:20], part_p[10][62]);
part_product p1063(move_ex[10][63:62], Y[22:20], part_p[10][63]);
part_product p1064(move_ex[10][64:63], Y[22:20], part_p[10][64]);
part_product p1065(move_ex[10][65:64], Y[22:20], part_p[10][65]);
part_product p1066(move_ex[10][66:65], Y[22:20], part_p[10][66]);
part_product p1067(move_ex[10][67:66], Y[22:20], part_p[10][67]);
get_c getc10(Y[22:20], C[21:20]);

assign part_p[11][0] = 0;
assign part_p[11][1] = 0;
assign part_p[11][2] = 0;
assign part_p[11][3] = 0;
assign part_p[11][4] = 0;
assign part_p[11][5] = 0;
assign part_p[11][6] = 0;
assign part_p[11][7] = 0;
assign part_p[11][8] = 0;
assign part_p[11][9] = 0;
assign part_p[11][10] = 0;
assign part_p[11][11] = 0;
assign part_p[11][12] = 0;
assign part_p[11][13] = 0;
assign part_p[11][14] = 0;
assign part_p[11][15] = 0;
assign part_p[11][16] = 0;
assign part_p[11][17] = 0;
assign part_p[11][18] = 0;
assign part_p[11][19] = 0;
assign part_p[11][20] = 0;
assign part_p[11][21] = 0;
s_part_product sp1122(move_ex[11][22:22], Y[24:22], part_p[11][22]);
part_product p1123(move_ex[11][23:22], Y[24:22], part_p[11][23]);
part_product p1124(move_ex[11][24:23], Y[24:22], part_p[11][24]);
part_product p1125(move_ex[11][25:24], Y[24:22], part_p[11][25]);
part_product p1126(move_ex[11][26:25], Y[24:22], part_p[11][26]);
part_product p1127(move_ex[11][27:26], Y[24:22], part_p[11][27]);
part_product p1128(move_ex[11][28:27], Y[24:22], part_p[11][28]);
part_product p1129(move_ex[11][29:28], Y[24:22], part_p[11][29]);
part_product p1130(move_ex[11][30:29], Y[24:22], part_p[11][30]);
part_product p1131(move_ex[11][31:30], Y[24:22], part_p[11][31]);
part_product p1132(move_ex[11][32:31], Y[24:22], part_p[11][32]);
part_product p1133(move_ex[11][33:32], Y[24:22], part_p[11][33]);
part_product p1134(move_ex[11][34:33], Y[24:22], part_p[11][34]);
part_product p1135(move_ex[11][35:34], Y[24:22], part_p[11][35]);
part_product p1136(move_ex[11][36:35], Y[24:22], part_p[11][36]);
part_product p1137(move_ex[11][37:36], Y[24:22], part_p[11][37]);
part_product p1138(move_ex[11][38:37], Y[24:22], part_p[11][38]);
part_product p1139(move_ex[11][39:38], Y[24:22], part_p[11][39]);
part_product p1140(move_ex[11][40:39], Y[24:22], part_p[11][40]);
part_product p1141(move_ex[11][41:40], Y[24:22], part_p[11][41]);
part_product p1142(move_ex[11][42:41], Y[24:22], part_p[11][42]);
part_product p1143(move_ex[11][43:42], Y[24:22], part_p[11][43]);
part_product p1144(move_ex[11][44:43], Y[24:22], part_p[11][44]);
part_product p1145(move_ex[11][45:44], Y[24:22], part_p[11][45]);
part_product p1146(move_ex[11][46:45], Y[24:22], part_p[11][46]);
part_product p1147(move_ex[11][47:46], Y[24:22], part_p[11][47]);
part_product p1148(move_ex[11][48:47], Y[24:22], part_p[11][48]);
part_product p1149(move_ex[11][49:48], Y[24:22], part_p[11][49]);
part_product p1150(move_ex[11][50:49], Y[24:22], part_p[11][50]);
part_product p1151(move_ex[11][51:50], Y[24:22], part_p[11][51]);
part_product p1152(move_ex[11][52:51], Y[24:22], part_p[11][52]);
part_product p1153(move_ex[11][53:52], Y[24:22], part_p[11][53]);
part_product p1154(move_ex[11][54:53], Y[24:22], part_p[11][54]);
part_product p1155(move_ex[11][55:54], Y[24:22], part_p[11][55]);
part_product p1156(move_ex[11][56:55], Y[24:22], part_p[11][56]);
part_product p1157(move_ex[11][57:56], Y[24:22], part_p[11][57]);
part_product p1158(move_ex[11][58:57], Y[24:22], part_p[11][58]);
part_product p1159(move_ex[11][59:58], Y[24:22], part_p[11][59]);
part_product p1160(move_ex[11][60:59], Y[24:22], part_p[11][60]);
part_product p1161(move_ex[11][61:60], Y[24:22], part_p[11][61]);
part_product p1162(move_ex[11][62:61], Y[24:22], part_p[11][62]);
part_product p1163(move_ex[11][63:62], Y[24:22], part_p[11][63]);
part_product p1164(move_ex[11][64:63], Y[24:22], part_p[11][64]);
part_product p1165(move_ex[11][65:64], Y[24:22], part_p[11][65]);
part_product p1166(move_ex[11][66:65], Y[24:22], part_p[11][66]);
part_product p1167(move_ex[11][67:66], Y[24:22], part_p[11][67]);
get_c getc11(Y[24:22], C[23:22]);

assign part_p[12][0] = 0;
assign part_p[12][1] = 0;
assign part_p[12][2] = 0;
assign part_p[12][3] = 0;
assign part_p[12][4] = 0;
assign part_p[12][5] = 0;
assign part_p[12][6] = 0;
assign part_p[12][7] = 0;
assign part_p[12][8] = 0;
assign part_p[12][9] = 0;
assign part_p[12][10] = 0;
assign part_p[12][11] = 0;
assign part_p[12][12] = 0;
assign part_p[12][13] = 0;
assign part_p[12][14] = 0;
assign part_p[12][15] = 0;
assign part_p[12][16] = 0;
assign part_p[12][17] = 0;
assign part_p[12][18] = 0;
assign part_p[12][19] = 0;
assign part_p[12][20] = 0;
assign part_p[12][21] = 0;
assign part_p[12][22] = 0;
assign part_p[12][23] = 0;
s_part_product sp1224(move_ex[12][24:24], Y[26:24], part_p[12][24]);
part_product p1225(move_ex[12][25:24], Y[26:24], part_p[12][25]);
part_product p1226(move_ex[12][26:25], Y[26:24], part_p[12][26]);
part_product p1227(move_ex[12][27:26], Y[26:24], part_p[12][27]);
part_product p1228(move_ex[12][28:27], Y[26:24], part_p[12][28]);
part_product p1229(move_ex[12][29:28], Y[26:24], part_p[12][29]);
part_product p1230(move_ex[12][30:29], Y[26:24], part_p[12][30]);
part_product p1231(move_ex[12][31:30], Y[26:24], part_p[12][31]);
part_product p1232(move_ex[12][32:31], Y[26:24], part_p[12][32]);
part_product p1233(move_ex[12][33:32], Y[26:24], part_p[12][33]);
part_product p1234(move_ex[12][34:33], Y[26:24], part_p[12][34]);
part_product p1235(move_ex[12][35:34], Y[26:24], part_p[12][35]);
part_product p1236(move_ex[12][36:35], Y[26:24], part_p[12][36]);
part_product p1237(move_ex[12][37:36], Y[26:24], part_p[12][37]);
part_product p1238(move_ex[12][38:37], Y[26:24], part_p[12][38]);
part_product p1239(move_ex[12][39:38], Y[26:24], part_p[12][39]);
part_product p1240(move_ex[12][40:39], Y[26:24], part_p[12][40]);
part_product p1241(move_ex[12][41:40], Y[26:24], part_p[12][41]);
part_product p1242(move_ex[12][42:41], Y[26:24], part_p[12][42]);
part_product p1243(move_ex[12][43:42], Y[26:24], part_p[12][43]);
part_product p1244(move_ex[12][44:43], Y[26:24], part_p[12][44]);
part_product p1245(move_ex[12][45:44], Y[26:24], part_p[12][45]);
part_product p1246(move_ex[12][46:45], Y[26:24], part_p[12][46]);
part_product p1247(move_ex[12][47:46], Y[26:24], part_p[12][47]);
part_product p1248(move_ex[12][48:47], Y[26:24], part_p[12][48]);
part_product p1249(move_ex[12][49:48], Y[26:24], part_p[12][49]);
part_product p1250(move_ex[12][50:49], Y[26:24], part_p[12][50]);
part_product p1251(move_ex[12][51:50], Y[26:24], part_p[12][51]);
part_product p1252(move_ex[12][52:51], Y[26:24], part_p[12][52]);
part_product p1253(move_ex[12][53:52], Y[26:24], part_p[12][53]);
part_product p1254(move_ex[12][54:53], Y[26:24], part_p[12][54]);
part_product p1255(move_ex[12][55:54], Y[26:24], part_p[12][55]);
part_product p1256(move_ex[12][56:55], Y[26:24], part_p[12][56]);
part_product p1257(move_ex[12][57:56], Y[26:24], part_p[12][57]);
part_product p1258(move_ex[12][58:57], Y[26:24], part_p[12][58]);
part_product p1259(move_ex[12][59:58], Y[26:24], part_p[12][59]);
part_product p1260(move_ex[12][60:59], Y[26:24], part_p[12][60]);
part_product p1261(move_ex[12][61:60], Y[26:24], part_p[12][61]);
part_product p1262(move_ex[12][62:61], Y[26:24], part_p[12][62]);
part_product p1263(move_ex[12][63:62], Y[26:24], part_p[12][63]);
part_product p1264(move_ex[12][64:63], Y[26:24], part_p[12][64]);
part_product p1265(move_ex[12][65:64], Y[26:24], part_p[12][65]);
part_product p1266(move_ex[12][66:65], Y[26:24], part_p[12][66]);
part_product p1267(move_ex[12][67:66], Y[26:24], part_p[12][67]);
get_c getc12(Y[26:24], C[25:24]);

assign part_p[13][0] = 0;
assign part_p[13][1] = 0;
assign part_p[13][2] = 0;
assign part_p[13][3] = 0;
assign part_p[13][4] = 0;
assign part_p[13][5] = 0;
assign part_p[13][6] = 0;
assign part_p[13][7] = 0;
assign part_p[13][8] = 0;
assign part_p[13][9] = 0;
assign part_p[13][10] = 0;
assign part_p[13][11] = 0;
assign part_p[13][12] = 0;
assign part_p[13][13] = 0;
assign part_p[13][14] = 0;
assign part_p[13][15] = 0;
assign part_p[13][16] = 0;
assign part_p[13][17] = 0;
assign part_p[13][18] = 0;
assign part_p[13][19] = 0;
assign part_p[13][20] = 0;
assign part_p[13][21] = 0;
assign part_p[13][22] = 0;
assign part_p[13][23] = 0;
assign part_p[13][24] = 0;
assign part_p[13][25] = 0;
s_part_product sp1326(move_ex[13][26:26], Y[28:26], part_p[13][26]);
part_product p1327(move_ex[13][27:26], Y[28:26], part_p[13][27]);
part_product p1328(move_ex[13][28:27], Y[28:26], part_p[13][28]);
part_product p1329(move_ex[13][29:28], Y[28:26], part_p[13][29]);
part_product p1330(move_ex[13][30:29], Y[28:26], part_p[13][30]);
part_product p1331(move_ex[13][31:30], Y[28:26], part_p[13][31]);
part_product p1332(move_ex[13][32:31], Y[28:26], part_p[13][32]);
part_product p1333(move_ex[13][33:32], Y[28:26], part_p[13][33]);
part_product p1334(move_ex[13][34:33], Y[28:26], part_p[13][34]);
part_product p1335(move_ex[13][35:34], Y[28:26], part_p[13][35]);
part_product p1336(move_ex[13][36:35], Y[28:26], part_p[13][36]);
part_product p1337(move_ex[13][37:36], Y[28:26], part_p[13][37]);
part_product p1338(move_ex[13][38:37], Y[28:26], part_p[13][38]);
part_product p1339(move_ex[13][39:38], Y[28:26], part_p[13][39]);
part_product p1340(move_ex[13][40:39], Y[28:26], part_p[13][40]);
part_product p1341(move_ex[13][41:40], Y[28:26], part_p[13][41]);
part_product p1342(move_ex[13][42:41], Y[28:26], part_p[13][42]);
part_product p1343(move_ex[13][43:42], Y[28:26], part_p[13][43]);
part_product p1344(move_ex[13][44:43], Y[28:26], part_p[13][44]);
part_product p1345(move_ex[13][45:44], Y[28:26], part_p[13][45]);
part_product p1346(move_ex[13][46:45], Y[28:26], part_p[13][46]);
part_product p1347(move_ex[13][47:46], Y[28:26], part_p[13][47]);
part_product p1348(move_ex[13][48:47], Y[28:26], part_p[13][48]);
part_product p1349(move_ex[13][49:48], Y[28:26], part_p[13][49]);
part_product p1350(move_ex[13][50:49], Y[28:26], part_p[13][50]);
part_product p1351(move_ex[13][51:50], Y[28:26], part_p[13][51]);
part_product p1352(move_ex[13][52:51], Y[28:26], part_p[13][52]);
part_product p1353(move_ex[13][53:52], Y[28:26], part_p[13][53]);
part_product p1354(move_ex[13][54:53], Y[28:26], part_p[13][54]);
part_product p1355(move_ex[13][55:54], Y[28:26], part_p[13][55]);
part_product p1356(move_ex[13][56:55], Y[28:26], part_p[13][56]);
part_product p1357(move_ex[13][57:56], Y[28:26], part_p[13][57]);
part_product p1358(move_ex[13][58:57], Y[28:26], part_p[13][58]);
part_product p1359(move_ex[13][59:58], Y[28:26], part_p[13][59]);
part_product p1360(move_ex[13][60:59], Y[28:26], part_p[13][60]);
part_product p1361(move_ex[13][61:60], Y[28:26], part_p[13][61]);
part_product p1362(move_ex[13][62:61], Y[28:26], part_p[13][62]);
part_product p1363(move_ex[13][63:62], Y[28:26], part_p[13][63]);
part_product p1364(move_ex[13][64:63], Y[28:26], part_p[13][64]);
part_product p1365(move_ex[13][65:64], Y[28:26], part_p[13][65]);
part_product p1366(move_ex[13][66:65], Y[28:26], part_p[13][66]);
part_product p1367(move_ex[13][67:66], Y[28:26], part_p[13][67]);
get_c getc13(Y[28:26], C[27:26]);

assign part_p[14][0] = 0;
assign part_p[14][1] = 0;
assign part_p[14][2] = 0;
assign part_p[14][3] = 0;
assign part_p[14][4] = 0;
assign part_p[14][5] = 0;
assign part_p[14][6] = 0;
assign part_p[14][7] = 0;
assign part_p[14][8] = 0;
assign part_p[14][9] = 0;
assign part_p[14][10] = 0;
assign part_p[14][11] = 0;
assign part_p[14][12] = 0;
assign part_p[14][13] = 0;
assign part_p[14][14] = 0;
assign part_p[14][15] = 0;
assign part_p[14][16] = 0;
assign part_p[14][17] = 0;
assign part_p[14][18] = 0;
assign part_p[14][19] = 0;
assign part_p[14][20] = 0;
assign part_p[14][21] = 0;
assign part_p[14][22] = 0;
assign part_p[14][23] = 0;
assign part_p[14][24] = 0;
assign part_p[14][25] = 0;
assign part_p[14][26] = 0;
assign part_p[14][27] = 0;
s_part_product sp1428(move_ex[14][28:28], Y[30:28], part_p[14][28]);
part_product p1429(move_ex[14][29:28], Y[30:28], part_p[14][29]);
part_product p1430(move_ex[14][30:29], Y[30:28], part_p[14][30]);
part_product p1431(move_ex[14][31:30], Y[30:28], part_p[14][31]);
part_product p1432(move_ex[14][32:31], Y[30:28], part_p[14][32]);
part_product p1433(move_ex[14][33:32], Y[30:28], part_p[14][33]);
part_product p1434(move_ex[14][34:33], Y[30:28], part_p[14][34]);
part_product p1435(move_ex[14][35:34], Y[30:28], part_p[14][35]);
part_product p1436(move_ex[14][36:35], Y[30:28], part_p[14][36]);
part_product p1437(move_ex[14][37:36], Y[30:28], part_p[14][37]);
part_product p1438(move_ex[14][38:37], Y[30:28], part_p[14][38]);
part_product p1439(move_ex[14][39:38], Y[30:28], part_p[14][39]);
part_product p1440(move_ex[14][40:39], Y[30:28], part_p[14][40]);
part_product p1441(move_ex[14][41:40], Y[30:28], part_p[14][41]);
part_product p1442(move_ex[14][42:41], Y[30:28], part_p[14][42]);
part_product p1443(move_ex[14][43:42], Y[30:28], part_p[14][43]);
part_product p1444(move_ex[14][44:43], Y[30:28], part_p[14][44]);
part_product p1445(move_ex[14][45:44], Y[30:28], part_p[14][45]);
part_product p1446(move_ex[14][46:45], Y[30:28], part_p[14][46]);
part_product p1447(move_ex[14][47:46], Y[30:28], part_p[14][47]);
part_product p1448(move_ex[14][48:47], Y[30:28], part_p[14][48]);
part_product p1449(move_ex[14][49:48], Y[30:28], part_p[14][49]);
part_product p1450(move_ex[14][50:49], Y[30:28], part_p[14][50]);
part_product p1451(move_ex[14][51:50], Y[30:28], part_p[14][51]);
part_product p1452(move_ex[14][52:51], Y[30:28], part_p[14][52]);
part_product p1453(move_ex[14][53:52], Y[30:28], part_p[14][53]);
part_product p1454(move_ex[14][54:53], Y[30:28], part_p[14][54]);
part_product p1455(move_ex[14][55:54], Y[30:28], part_p[14][55]);
part_product p1456(move_ex[14][56:55], Y[30:28], part_p[14][56]);
part_product p1457(move_ex[14][57:56], Y[30:28], part_p[14][57]);
part_product p1458(move_ex[14][58:57], Y[30:28], part_p[14][58]);
part_product p1459(move_ex[14][59:58], Y[30:28], part_p[14][59]);
part_product p1460(move_ex[14][60:59], Y[30:28], part_p[14][60]);
part_product p1461(move_ex[14][61:60], Y[30:28], part_p[14][61]);
part_product p1462(move_ex[14][62:61], Y[30:28], part_p[14][62]);
part_product p1463(move_ex[14][63:62], Y[30:28], part_p[14][63]);
part_product p1464(move_ex[14][64:63], Y[30:28], part_p[14][64]);
part_product p1465(move_ex[14][65:64], Y[30:28], part_p[14][65]);
part_product p1466(move_ex[14][66:65], Y[30:28], part_p[14][66]);
part_product p1467(move_ex[14][67:66], Y[30:28], part_p[14][67]);
get_c getc14(Y[30:28], C[29:28]);

assign part_p[15][0] = 0;
assign part_p[15][1] = 0;
assign part_p[15][2] = 0;
assign part_p[15][3] = 0;
assign part_p[15][4] = 0;
assign part_p[15][5] = 0;
assign part_p[15][6] = 0;
assign part_p[15][7] = 0;
assign part_p[15][8] = 0;
assign part_p[15][9] = 0;
assign part_p[15][10] = 0;
assign part_p[15][11] = 0;
assign part_p[15][12] = 0;
assign part_p[15][13] = 0;
assign part_p[15][14] = 0;
assign part_p[15][15] = 0;
assign part_p[15][16] = 0;
assign part_p[15][17] = 0;
assign part_p[15][18] = 0;
assign part_p[15][19] = 0;
assign part_p[15][20] = 0;
assign part_p[15][21] = 0;
assign part_p[15][22] = 0;
assign part_p[15][23] = 0;
assign part_p[15][24] = 0;
assign part_p[15][25] = 0;
assign part_p[15][26] = 0;
assign part_p[15][27] = 0;
assign part_p[15][28] = 0;
assign part_p[15][29] = 0;
s_part_product sp1530(move_ex[15][30:30], Y[32:30], part_p[15][30]);
part_product p1531(move_ex[15][31:30], Y[32:30], part_p[15][31]);
part_product p1532(move_ex[15][32:31], Y[32:30], part_p[15][32]);
part_product p1533(move_ex[15][33:32], Y[32:30], part_p[15][33]);
part_product p1534(move_ex[15][34:33], Y[32:30], part_p[15][34]);
part_product p1535(move_ex[15][35:34], Y[32:30], part_p[15][35]);
part_product p1536(move_ex[15][36:35], Y[32:30], part_p[15][36]);
part_product p1537(move_ex[15][37:36], Y[32:30], part_p[15][37]);
part_product p1538(move_ex[15][38:37], Y[32:30], part_p[15][38]);
part_product p1539(move_ex[15][39:38], Y[32:30], part_p[15][39]);
part_product p1540(move_ex[15][40:39], Y[32:30], part_p[15][40]);
part_product p1541(move_ex[15][41:40], Y[32:30], part_p[15][41]);
part_product p1542(move_ex[15][42:41], Y[32:30], part_p[15][42]);
part_product p1543(move_ex[15][43:42], Y[32:30], part_p[15][43]);
part_product p1544(move_ex[15][44:43], Y[32:30], part_p[15][44]);
part_product p1545(move_ex[15][45:44], Y[32:30], part_p[15][45]);
part_product p1546(move_ex[15][46:45], Y[32:30], part_p[15][46]);
part_product p1547(move_ex[15][47:46], Y[32:30], part_p[15][47]);
part_product p1548(move_ex[15][48:47], Y[32:30], part_p[15][48]);
part_product p1549(move_ex[15][49:48], Y[32:30], part_p[15][49]);
part_product p1550(move_ex[15][50:49], Y[32:30], part_p[15][50]);
part_product p1551(move_ex[15][51:50], Y[32:30], part_p[15][51]);
part_product p1552(move_ex[15][52:51], Y[32:30], part_p[15][52]);
part_product p1553(move_ex[15][53:52], Y[32:30], part_p[15][53]);
part_product p1554(move_ex[15][54:53], Y[32:30], part_p[15][54]);
part_product p1555(move_ex[15][55:54], Y[32:30], part_p[15][55]);
part_product p1556(move_ex[15][56:55], Y[32:30], part_p[15][56]);
part_product p1557(move_ex[15][57:56], Y[32:30], part_p[15][57]);
part_product p1558(move_ex[15][58:57], Y[32:30], part_p[15][58]);
part_product p1559(move_ex[15][59:58], Y[32:30], part_p[15][59]);
part_product p1560(move_ex[15][60:59], Y[32:30], part_p[15][60]);
part_product p1561(move_ex[15][61:60], Y[32:30], part_p[15][61]);
part_product p1562(move_ex[15][62:61], Y[32:30], part_p[15][62]);
part_product p1563(move_ex[15][63:62], Y[32:30], part_p[15][63]);
part_product p1564(move_ex[15][64:63], Y[32:30], part_p[15][64]);
part_product p1565(move_ex[15][65:64], Y[32:30], part_p[15][65]);
part_product p1566(move_ex[15][66:65], Y[32:30], part_p[15][66]);
part_product p1567(move_ex[15][67:66], Y[32:30], part_p[15][67]);
get_c getc15(Y[32:30], C[31:30]);

assign part_p[16][0] = 0;
assign part_p[16][1] = 0;
assign part_p[16][2] = 0;
assign part_p[16][3] = 0;
assign part_p[16][4] = 0;
assign part_p[16][5] = 0;
assign part_p[16][6] = 0;
assign part_p[16][7] = 0;
assign part_p[16][8] = 0;
assign part_p[16][9] = 0;
assign part_p[16][10] = 0;
assign part_p[16][11] = 0;
assign part_p[16][12] = 0;
assign part_p[16][13] = 0;
assign part_p[16][14] = 0;
assign part_p[16][15] = 0;
assign part_p[16][16] = 0;
assign part_p[16][17] = 0;
assign part_p[16][18] = 0;
assign part_p[16][19] = 0;
assign part_p[16][20] = 0;
assign part_p[16][21] = 0;
assign part_p[16][22] = 0;
assign part_p[16][23] = 0;
assign part_p[16][24] = 0;
assign part_p[16][25] = 0;
assign part_p[16][26] = 0;
assign part_p[16][27] = 0;
assign part_p[16][28] = 0;
assign part_p[16][29] = 0;
assign part_p[16][30] = 0;
assign part_p[16][31] = 0;
s_part_product sp1632(move_ex[16][32:32], Y[34:32], part_p[16][32]);
part_product p1633(move_ex[16][33:32], Y[34:32], part_p[16][33]);
part_product p1634(move_ex[16][34:33], Y[34:32], part_p[16][34]);
part_product p1635(move_ex[16][35:34], Y[34:32], part_p[16][35]);
part_product p1636(move_ex[16][36:35], Y[34:32], part_p[16][36]);
part_product p1637(move_ex[16][37:36], Y[34:32], part_p[16][37]);
part_product p1638(move_ex[16][38:37], Y[34:32], part_p[16][38]);
part_product p1639(move_ex[16][39:38], Y[34:32], part_p[16][39]);
part_product p1640(move_ex[16][40:39], Y[34:32], part_p[16][40]);
part_product p1641(move_ex[16][41:40], Y[34:32], part_p[16][41]);
part_product p1642(move_ex[16][42:41], Y[34:32], part_p[16][42]);
part_product p1643(move_ex[16][43:42], Y[34:32], part_p[16][43]);
part_product p1644(move_ex[16][44:43], Y[34:32], part_p[16][44]);
part_product p1645(move_ex[16][45:44], Y[34:32], part_p[16][45]);
part_product p1646(move_ex[16][46:45], Y[34:32], part_p[16][46]);
part_product p1647(move_ex[16][47:46], Y[34:32], part_p[16][47]);
part_product p1648(move_ex[16][48:47], Y[34:32], part_p[16][48]);
part_product p1649(move_ex[16][49:48], Y[34:32], part_p[16][49]);
part_product p1650(move_ex[16][50:49], Y[34:32], part_p[16][50]);
part_product p1651(move_ex[16][51:50], Y[34:32], part_p[16][51]);
part_product p1652(move_ex[16][52:51], Y[34:32], part_p[16][52]);
part_product p1653(move_ex[16][53:52], Y[34:32], part_p[16][53]);
part_product p1654(move_ex[16][54:53], Y[34:32], part_p[16][54]);
part_product p1655(move_ex[16][55:54], Y[34:32], part_p[16][55]);
part_product p1656(move_ex[16][56:55], Y[34:32], part_p[16][56]);
part_product p1657(move_ex[16][57:56], Y[34:32], part_p[16][57]);
part_product p1658(move_ex[16][58:57], Y[34:32], part_p[16][58]);
part_product p1659(move_ex[16][59:58], Y[34:32], part_p[16][59]);
part_product p1660(move_ex[16][60:59], Y[34:32], part_p[16][60]);
part_product p1661(move_ex[16][61:60], Y[34:32], part_p[16][61]);
part_product p1662(move_ex[16][62:61], Y[34:32], part_p[16][62]);
part_product p1663(move_ex[16][63:62], Y[34:32], part_p[16][63]);
part_product p1664(move_ex[16][64:63], Y[34:32], part_p[16][64]);
part_product p1665(move_ex[16][65:64], Y[34:32], part_p[16][65]);
part_product p1666(move_ex[16][66:65], Y[34:32], part_p[16][66]);
part_product p1667(move_ex[16][67:66], Y[34:32], part_p[16][67]);
get_c getc16(Y[34:32], C[33:32]);
assign C[67:34] = 0;




wire [16:0] new_p[0:67];
switch sw(part_p[0], part_p[1], part_p[2], part_p[3], part_p[4], part_p[5], part_p[6], part_p[7], part_p[8], part_p[9], part_p[10], part_p[11], part_p[12], part_p[13], part_p[14], part_p[15], part_p[16], new_p[0], new_p[1], new_p[2], new_p[3], new_p[4], new_p[5], new_p[6], new_p[7], new_p[8], new_p[9], new_p[10], new_p[11], new_p[12], new_p[13], new_p[14], new_p[15], new_p[16], new_p[17], new_p[18], new_p[19], new_p[20], new_p[21], new_p[22], new_p[23], new_p[24], new_p[25], new_p[26], new_p[27], new_p[28], new_p[29], new_p[30], new_p[31], new_p[32], new_p[33], new_p[34], new_p[35], new_p[36], new_p[37], new_p[38], new_p[39], new_p[40], new_p[41], new_p[42], new_p[43], new_p[44], new_p[45], new_p[46], new_p[47], new_p[48], new_p[49], new_p[50], new_p[51], new_p[52], new_p[53], new_p[54], new_p[55], new_p[56], new_p[57], new_p[58], new_p[59], new_p[60], new_p[61], new_p[62], new_p[63], new_p[64], new_p[65], new_p[66], new_p[67]);

wire [67:0] s, carry;
wire [13:0] cout [0:67];
walloc_17bits w17_0(new_p[0], 14'b0, cout[0], carry[0], s[0]);
walloc_17bits w17_1(new_p[1], cout[0], cout[1], carry[1], s[1]);
walloc_17bits w17_2(new_p[2], cout[1], cout[2], carry[2], s[2]);
walloc_17bits w17_3(new_p[3], cout[2], cout[3], carry[3], s[3]);
walloc_17bits w17_4(new_p[4], cout[3], cout[4], carry[4], s[4]);
walloc_17bits w17_5(new_p[5], cout[4], cout[5], carry[5], s[5]);
walloc_17bits w17_6(new_p[6], cout[5], cout[6], carry[6], s[6]);
walloc_17bits w17_7(new_p[7], cout[6], cout[7], carry[7], s[7]);
walloc_17bits w17_8(new_p[8], cout[7], cout[8], carry[8], s[8]);
walloc_17bits w17_9(new_p[9], cout[8], cout[9], carry[9], s[9]);
walloc_17bits w17_10(new_p[10], cout[9], cout[10], carry[10], s[10]);
walloc_17bits w17_11(new_p[11], cout[10], cout[11], carry[11], s[11]);
walloc_17bits w17_12(new_p[12], cout[11], cout[12], carry[12], s[12]);
walloc_17bits w17_13(new_p[13], cout[12], cout[13], carry[13], s[13]);
walloc_17bits w17_14(new_p[14], cout[13], cout[14], carry[14], s[14]);
walloc_17bits w17_15(new_p[15], cout[14], cout[15], carry[15], s[15]);
walloc_17bits w17_16(new_p[16], cout[15], cout[16], carry[16], s[16]);
walloc_17bits w17_17(new_p[17], cout[16], cout[17], carry[17], s[17]);
walloc_17bits w17_18(new_p[18], cout[17], cout[18], carry[18], s[18]);
walloc_17bits w17_19(new_p[19], cout[18], cout[19], carry[19], s[19]);
walloc_17bits w17_20(new_p[20], cout[19], cout[20], carry[20], s[20]);
walloc_17bits w17_21(new_p[21], cout[20], cout[21], carry[21], s[21]);
walloc_17bits w17_22(new_p[22], cout[21], cout[22], carry[22], s[22]);
walloc_17bits w17_23(new_p[23], cout[22], cout[23], carry[23], s[23]);
walloc_17bits w17_24(new_p[24], cout[23], cout[24], carry[24], s[24]);
walloc_17bits w17_25(new_p[25], cout[24], cout[25], carry[25], s[25]);
walloc_17bits w17_26(new_p[26], cout[25], cout[26], carry[26], s[26]);
walloc_17bits w17_27(new_p[27], cout[26], cout[27], carry[27], s[27]);
walloc_17bits w17_28(new_p[28], cout[27], cout[28], carry[28], s[28]);
walloc_17bits w17_29(new_p[29], cout[28], cout[29], carry[29], s[29]);
walloc_17bits w17_30(new_p[30], cout[29], cout[30], carry[30], s[30]);
walloc_17bits w17_31(new_p[31], cout[30], cout[31], carry[31], s[31]);
walloc_17bits w17_32(new_p[32], cout[31], cout[32], carry[32], s[32]);
walloc_17bits w17_33(new_p[33], cout[32], cout[33], carry[33], s[33]);
walloc_17bits w17_34(new_p[34], cout[33], cout[34], carry[34], s[34]);
walloc_17bits w17_35(new_p[35], cout[34], cout[35], carry[35], s[35]);
walloc_17bits w17_36(new_p[36], cout[35], cout[36], carry[36], s[36]);
walloc_17bits w17_37(new_p[37], cout[36], cout[37], carry[37], s[37]);
walloc_17bits w17_38(new_p[38], cout[37], cout[38], carry[38], s[38]);
walloc_17bits w17_39(new_p[39], cout[38], cout[39], carry[39], s[39]);
walloc_17bits w17_40(new_p[40], cout[39], cout[40], carry[40], s[40]);
walloc_17bits w17_41(new_p[41], cout[40], cout[41], carry[41], s[41]);
walloc_17bits w17_42(new_p[42], cout[41], cout[42], carry[42], s[42]);
walloc_17bits w17_43(new_p[43], cout[42], cout[43], carry[43], s[43]);
walloc_17bits w17_44(new_p[44], cout[43], cout[44], carry[44], s[44]);
walloc_17bits w17_45(new_p[45], cout[44], cout[45], carry[45], s[45]);
walloc_17bits w17_46(new_p[46], cout[45], cout[46], carry[46], s[46]);
walloc_17bits w17_47(new_p[47], cout[46], cout[47], carry[47], s[47]);
walloc_17bits w17_48(new_p[48], cout[47], cout[48], carry[48], s[48]);
walloc_17bits w17_49(new_p[49], cout[48], cout[49], carry[49], s[49]);
walloc_17bits w17_50(new_p[50], cout[49], cout[50], carry[50], s[50]);
walloc_17bits w17_51(new_p[51], cout[50], cout[51], carry[51], s[51]);
walloc_17bits w17_52(new_p[52], cout[51], cout[52], carry[52], s[52]);
walloc_17bits w17_53(new_p[53], cout[52], cout[53], carry[53], s[53]);
walloc_17bits w17_54(new_p[54], cout[53], cout[54], carry[54], s[54]);
walloc_17bits w17_55(new_p[55], cout[54], cout[55], carry[55], s[55]);
walloc_17bits w17_56(new_p[56], cout[55], cout[56], carry[56], s[56]);
walloc_17bits w17_57(new_p[57], cout[56], cout[57], carry[57], s[57]);
walloc_17bits w17_58(new_p[58], cout[57], cout[58], carry[58], s[58]);
walloc_17bits w17_59(new_p[59], cout[58], cout[59], carry[59], s[59]);
walloc_17bits w17_60(new_p[60], cout[59], cout[60], carry[60], s[60]);
walloc_17bits w17_61(new_p[61], cout[60], cout[61], carry[61], s[61]);
walloc_17bits w17_62(new_p[62], cout[61], cout[62], carry[62], s[62]);
walloc_17bits w17_63(new_p[63], cout[62], cout[63], carry[63], s[63]);
walloc_17bits w17_64(new_p[64], cout[63], cout[64], carry[64], s[64]);
walloc_17bits w17_65(new_p[65], cout[64], cout[65], carry[65], s[65]);
walloc_17bits w17_66(new_p[66], cout[65], cout[66], carry[66], s[66]);
walloc_17bits w17_67(new_p[67], cout[66], cout[67], carry[67], s[67]);



wire [67:0] temp, ttemp;
cla_68bits cla68_0(s[67:0], {carry[66:0], 1'b0}, 1'b0, temp[67:0]);
cla_68bits cla68_1(temp, C, 1'b0, ttemp);
assign res = ttemp[63:0];
endmodule